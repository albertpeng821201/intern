// (c) Copyright 2012-2016 PRO DESIGN Electronic GmbH.                     
// All rights reserved.                                                    
//                                                                         
// This file is owned and controlled by ProDesign and must be used solely  
// for design, simulation, implementation and creation of design files     
// limited to profpga systems or technologies. Use with non-profpga        
// systems or technologies is expressly prohibited and immediately         
// terminates your license.                                                
//                                                                         
// PRODESIGN IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY 
// FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR PRODESIGN SYSTEMS. BY  
// PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             
// IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, PRODESIGN IS   
// MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      
// CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       
// RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION. PRODESIGN EXPRESSLY     
// DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   
// IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          
// REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         
// INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   
// PARTICULAR PURPOSE.                                                     
//                                                                         
// ProDesign products are not intended for use in life support appliances, 
// devices, or systems. Use in such applications are expressly             
// prohibited.                                                             
//                                                                         
// This file was generated by profpga_brdgen version 6.02 
//   on Mon May 15 18:13:22 2017 

`ifndef PD_MUXDEMUX_PARAM_VH
`define PD_MUXDEMUX_PARAM_VH

`include "pd_muxdemux.vh"

// pd_muxdemux parameters which are common to all FPGA technologies
`define PD_MUXDEMUX_MUX_TYPE `PD_MUXDEMUX_MUX_TYPE_ASYNCMUXSYSSYNCCLK
`define PD_MUXDEMUX_SIM_MODE `PD_MUXDEMUX_SIM_MODE_PRODUCTION
`define PD_MUXDEMUX_MUX_FACTOR 4
`define PD_MUXDEMUX_WORD_COUNT 1
`define PD_MUXDEMUX_MIN_DATARATE_MBIT 600000000
`define PD_MUXDEMUX_MAX_DATARATE_MBIT 800000000
`define PD_MUXDEMUX_MIN_CLK_BASE_FREQUENCY_HZ 50000000
`define PD_MUXDEMUX_MAX_CLK_BASE_FREQUENCY_HZ 66666666
`define PD_MUXDEMUX_MIN_CLK_BASE_PERIOD_NS 20.000
`define PD_MUXDEMUX_MAX_CLK_BASE_PERIOD_NS 15.001

// dbst parameters
`define DBST_REVERSE_DIRECTION 0
`define DBST_IOSTANDARD 'h01 // SSTL18_I_DCI

// pd_muxdemux parameters which are dedicated to the FPGA module
//   MB_1.TA1
`define PD_MUXDEMUX_FPGA_TYPE "XC7V2000T"
`define PD_MUXDEMUX_FPGA_SPEED_GRADE 1
`define PD_MUXDEMUX_FPGA_TECHNOLOGY `PD_MUXDEMUX_FPGA_TECHNOLOGY_XV7

`define PD_MUXDEMUX_SERDES_MODE "DDR"
`define PD_MUXDEMUX_SERDES_MODE_BIT 1'b1
`define PD_MUXDEMUX_SERDES_FACTOR 4
`define PD_MUXDEMUX_PLL_M 24
`define PD_MUXDEMUX_PLL_D0 24
`define PD_MUXDEMUX_PLL_D1 4
`define PD_MUXDEMUX_PLL_D2 8
`define PD_MUXDEMUX_PLL_D3 24
`define PD_MUXDEMUX_ENABLE_DCIRESET 0

`endif
