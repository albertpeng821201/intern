/* (c) Copyright 2012-2016 PRO DESIGN Electronic GmbH.                     */
/* All rights reserved.                                                    */
/*                                                                         */
/* This file is owned and controlled by ProDesign and must be used solely  */
/* for design, simulation, implementation and creation of design files     */
/* limited to profpga systems or technologies. Use with non-profpga        */
/* systems or technologies is expressly prohibited and immediately         */
/* terminates your license.                                                */
/*                                                                         */
/* PRODESIGN IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY */
/* FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR PRODESIGN SYSTEMS. BY  */
/* PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             */
/* IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, PRODESIGN IS   */
/* MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      */
/* CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       */
/* RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION. PRODESIGN EXPRESSLY     */
/* DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   */
/* IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          */
/* REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         */
/* INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   */
/* PARTICULAR PURPOSE.                                                     */
/*                                                                         */
/* ProDesign products are not intended for use in life support appliances, */
/* devices, or systems. Use in such applications are expressly             */
/* prohibited.                                                             */
/*                                                                         */
/* This file was generated by profpga_brdgen version 6.02 */
/*   on Wed Mar 15 14:30:12 2017 */

import functions::*;
import types::*;
import parameters::*;

/* FPGA module FM-XC7V2000T-R2 */
module mb_1_TC3 (
    clk0_p,
    clk0_n,

    sync0_p,
    sync0_n,

    dmbi_h2f,
    dmbi_f2h,

    clk1_p,
    clk1_n,

    sync1_p,
    sync1_n,

    led_red,
    led_green,
    led_blue,
    led_yellow,

    `ifdef EN_DDR
        clk2_p,
        clk2_n,
    `endif

    // SSRAM interface
    sram0_k_p,
    sram0_k_n,
    sram0_a,
    sram0_dq,
    sram0_bws_n,
    sram0_rnw,
    sram0_ld_n,
    sram0_doff_n,

    sram1_k_p,
    sram1_k_n,
    sram1_a,
    sram1_dq,
    sram1_bws_n,
    sram1_rnw,
    sram1_ld_n,
    sram1_doff_n,

    sram2_k_p,
    sram2_k_n,
    sram2_a,
    sram2_dq,
    sram2_bws_n,
    sram2_rnw,
    sram2_ld_n,
    sram2_doff_n,

    sram3_k_p,
    sram3_k_n,
    sram3_a,
    sram3_dq,
    sram3_bws_n,
    sram3_rnw,
    sram3_ld_n,
    sram3_doff_n,

    `ifdef EN_DDR
        ddr3_dq,
        ddr3_dqs_p,
        ddr3_dqs_n,
        ddr3_addr,
        ddr3_ba ,
        ddr3_ras_n,
        ddr3_cas_n ,
        ddr3_we_n   ,
        ddr3_reset_n,
        ddr3_ck_p,
        ddr3_ck_n,
        ddr3_cke ,
        ddr3_cs_n ,
        ddr3_dm ,
        ddr3_odt,
    `endif

    `ifdef EN_ETH
        eth_clk_to_mac,
        eth_col_clk_mac_freq,
        eth_crs_rgmii_sel0,
        eth_gtx_clk_tck,
        eth_mdc,
        eth_mdio,
        eth_ninterrupt,
        eth_nreset,
        eth_rx_clk,
        eth_rx_dv_rck,
        eth_rx_er_rxdv_er,
        eth_rxd,
        eth_tx_clk_rgmii_sel1,
        eth_tx_en_txen_er,
        eth_tx_er,
        eth_txd,
    `endif

    mb1_BA3_CLKIO_N_0_mb1_BC3_CLKIO_N_7,  /* BA3_CLKIO_N_0 */
    mb1_BA3_CLKIO_N_1_mb1_BC3_CLKIO_N_6,  /* BA3_CLKIO_N_1 */
    mb1_BA3_CLKIO_N_2_mb1_BC3_CLKIO_N_4,  /* BA3_CLKIO_N_2 */
    mb1_BA3_CLKIO_N_3_mb1_BC3_CLKIO_N_3,  /* BA3_CLKIO_N_3 */
    mb1_BA3_CLKIO_N_4_mb1_BC3_CLKIO_N_2,  /* BA3_CLKIO_N_4 */
    mb1_BA3_CLKIO_N_5_mb1_BC3_IO_010,  /* BA3_CLKIO_N_5 */
    mb1_BA3_CLKIO_N_6_mb1_BC3_CLKIO_N_1,  /* BA3_CLKIO_N_6 */
    mb1_BA3_CLKIO_N_7_mb1_BC3_CLKIO_N_0,  /* BA3_CLKIO_N_7 */
    mb1_BA3_CLKIO_P_0_mb1_BC3_CLKIO_P_7,  /* BA3_CLKIO_P_0 */
    mb1_BA3_CLKIO_P_1_mb1_BC3_CLKIO_P_6,  /* BA3_CLKIO_P_1 */
    mb1_BA3_CLKIO_P_2_mb1_BC3_CLKIO_P_4,  /* BA3_CLKIO_P_2 */
    mb1_BA3_CLKIO_P_3_mb1_BC3_CLKIO_P_3,  /* BA3_CLKIO_P_3 */
    mb1_BA3_CLKIO_P_4_mb1_BC3_CLKIO_P_2,  /* BA3_CLKIO_P_4 */
    mb1_BA3_CLKIO_P_5_mb1_BC3_IO_011,  /* BA3_CLKIO_P_5 */
    mb1_BA3_CLKIO_P_6_mb1_BC3_CLKIO_P_1,  /* BA3_CLKIO_P_6 */
    mb1_BA3_CLKIO_P_7_mb1_BC3_CLKIO_P_0,  /* BA3_CLKIO_P_7 */
    mb1_BA3_IO_004_mb1_BC3_IO_006,  /* BA3_IO_004 */
    mb1_BA3_IO_005_mb1_BC3_IO_007,  /* BA3_IO_005 */
    mb1_BA3_IO_006_mb1_BC3_IO_004,  /* BA3_IO_006 */
    mb1_BA3_IO_007_mb1_BC3_IO_005,  /* BA3_IO_007 */
    mb1_BA3_IO_008_mb1_BC3_IO_022,  /* BA3_IO_008 */
    mb1_BA3_IO_009_mb1_BC3_IO_023,  /* BA3_IO_009 */
    mb1_BA3_IO_010_mb1_BC3_CLKIO_N_5,  /* BA3_IO_010 */
    mb1_BA3_IO_011_mb1_BC3_CLKIO_P_5,  /* BA3_IO_011 */
    mb1_BA3_IO_012_mb1_BC3_IO_012,  /* BA3_IO_012 */
    mb1_BA3_IO_013_mb1_BC3_IO_013,  /* BA3_IO_013 */
    mb1_BA3_IO_014_mb1_BC3_IO_016,  /* BA3_IO_014 */
    mb1_BA3_IO_015_mb1_BC3_IO_017,  /* BA3_IO_015 */
    mb1_BA3_IO_016_mb1_BC3_IO_014,  /* BA3_IO_016 */
    mb1_BA3_IO_017_mb1_BC3_IO_015,  /* BA3_IO_017 */
    mb1_BA3_IO_018_mb1_BC3_IO_032,  /* BA3_IO_018 */
    mb1_BA3_IO_019_mb1_BC3_IO_033,  /* BA3_IO_019 */
    mb1_BA3_IO_020_mb1_BC3_IO_030,  /* BA3_IO_020 */
    mb1_BA3_IO_021_mb1_BC3_IO_031,  /* BA3_IO_021 */
    mb1_BA3_IO_022_mb1_BC3_IO_008,  /* BA3_IO_022 */
    mb1_BA3_IO_023_mb1_BC3_IO_009,  /* BA3_IO_023 */
    mb1_BA3_IO_024_mb1_BC3_IO_026,  /* BA3_IO_024 */
    mb1_BA3_IO_025_mb1_BC3_IO_027,  /* BA3_IO_025 */
    mb1_BA3_IO_026_mb1_BC3_IO_024,  /* BA3_IO_026 */
    mb1_BA3_IO_027_mb1_BC3_IO_025,  /* BA3_IO_027 */
    mb1_BA3_IO_028_mb1_BC3_IO_042,  /* BA3_IO_028 */
    mb1_BA3_IO_029_mb1_BC3_IO_043,  /* BA3_IO_029 */
    mb1_BA3_IO_030_mb1_BC3_IO_020,  /* BA3_IO_030 */
    mb1_BA3_IO_031_mb1_BC3_IO_021,  /* BA3_IO_031 */
    mb1_BA3_IO_032_mb1_BC3_IO_018,  /* BA3_IO_032 */
    mb1_BA3_IO_033_mb1_BC3_IO_019,  /* BA3_IO_033 */
    mb1_BA3_IO_034_mb1_BC3_IO_036,  /* BA3_IO_034 */
    mb1_BA3_IO_035_mb1_BC3_IO_037,  /* BA3_IO_035 */
    mb1_BA3_IO_036_mb1_BC3_IO_034,  /* BA3_IO_036 */
    mb1_BA3_IO_037_mb1_BC3_IO_035,  /* BA3_IO_037 */
    mb1_BA3_IO_038_mb1_BC3_IO_052,  /* BA3_IO_038 */
    mb1_BA3_IO_039_mb1_BC3_IO_053,  /* BA3_IO_039 */
    mb1_BA3_IO_040_mb1_BC3_IO_050,  /* BA3_IO_040 */
    mb1_BA3_IO_041_mb1_BC3_IO_051,  /* BA3_IO_041 */
    mb1_BA3_IO_042_mb1_BC3_IO_028,  /* BA3_IO_042 */
    mb1_BA3_IO_043_mb1_BC3_IO_029,  /* BA3_IO_043 */
    mb1_BA3_IO_044_mb1_BC3_IO_046,  /* BA3_IO_044 */
    mb1_BA3_IO_045_mb1_BC3_IO_047,  /* BA3_IO_045 */
    mb1_BA3_IO_046_mb1_BC3_IO_044,  /* BA3_IO_046 */
    mb1_BA3_IO_047_mb1_BC3_IO_045,  /* BA3_IO_047 */
    mb1_BA3_IO_048_mb1_BC3_IO_062,  /* BA3_IO_048 */
    mb1_BA3_IO_049_mb1_BC3_IO_063,  /* BA3_IO_049 */
    mb1_BA3_IO_050_mb1_BC3_IO_040,  /* BA3_IO_050 */
    mb1_BA3_IO_051_mb1_BC3_IO_041,  /* BA3_IO_051 */
    mb1_BA3_IO_052_mb1_BC3_IO_038,  /* BA3_IO_052 */
    mb1_BA3_IO_053_mb1_BC3_IO_039,  /* BA3_IO_053 */
    mb1_BA3_IO_054_mb1_BC3_IO_056,  /* BA3_IO_054 */
    mb1_BA3_IO_055_mb1_BC3_IO_057,  /* BA3_IO_055 */
    mb1_BA3_IO_056_mb1_BC3_IO_054,  /* BA3_IO_056 */
    mb1_BA3_IO_057_mb1_BC3_IO_055,  /* BA3_IO_057 */
    mb1_BA3_IO_058_mb1_BC3_IO_072,  /* BA3_IO_058 */
    mb1_BA3_IO_059_mb1_BC3_IO_073,  /* BA3_IO_059 */
    mb1_BA3_IO_060_mb1_BC3_IO_070,  /* BA3_IO_060 */
    mb1_BA3_IO_061_mb1_BC3_IO_071,  /* BA3_IO_061 */
    mb1_BA3_IO_062_mb1_BC3_IO_048,  /* BA3_IO_062 */
    mb1_BA3_IO_063_mb1_BC3_IO_049,  /* BA3_IO_063 */
    mb1_BA3_IO_064_mb1_BC3_IO_066,  /* BA3_IO_064 */
    mb1_BA3_IO_065_mb1_BC3_IO_067,  /* BA3_IO_065 */
    mb1_BA3_IO_066_mb1_BC3_IO_064,  /* BA3_IO_066 */
    mb1_BA3_IO_067_mb1_BC3_IO_065,  /* BA3_IO_067 */
    mb1_BA3_IO_068_mb1_BC3_IO_082,  /* BA3_IO_068 */
    mb1_BA3_IO_069_mb1_BC3_IO_083,  /* BA3_IO_069 */
    mb1_BA3_IO_070_mb1_BC3_IO_060,  /* BA3_IO_070 */
    mb1_BA3_IO_071_mb1_BC3_IO_061,  /* BA3_IO_071 */
    mb1_BA3_IO_072_mb1_BC3_IO_058,  /* BA3_IO_072 */
    mb1_BA3_IO_073_mb1_BC3_IO_059,  /* BA3_IO_073 */
    mb1_BA3_IO_074_mb1_BC3_IO_076,  /* BA3_IO_074 */
    mb1_BA3_IO_075_mb1_BC3_IO_077,  /* BA3_IO_075 */
    mb1_BA3_IO_076_mb1_BC3_IO_074,  /* BA3_IO_076 */
    mb1_BA3_IO_077_mb1_BC3_IO_075,  /* BA3_IO_077 */
    mb1_BA3_IO_078_mb1_BC3_IO_092,  /* BA3_IO_078 */
    mb1_BA3_IO_079_mb1_BC3_IO_093,  /* BA3_IO_079 */
    mb1_BA3_IO_080_mb1_BC3_IO_090,  /* BA3_IO_080 */
    mb1_BA3_IO_081_mb1_BC3_IO_091,  /* BA3_IO_081 */
    mb1_BA3_IO_082_mb1_BC3_IO_068,  /* BA3_IO_082 */
    mb1_BA3_IO_083_mb1_BC3_IO_069,  /* BA3_IO_083 */
    mb1_BA3_IO_084_mb1_BC3_IO_086,  /* BA3_IO_084 */
    mb1_BA3_IO_085_mb1_BC3_IO_087,  /* BA3_IO_085 */
    mb1_BA3_IO_086_mb1_BC3_IO_084,  /* BA3_IO_086 */
    mb1_BA3_IO_087_mb1_BC3_IO_085,  /* BA3_IO_087 */
    mb1_BA3_IO_088_mb1_BC3_IO_102,  /* BA3_IO_088 */
    mb1_BA3_IO_089_mb1_BC3_IO_103,  /* BA3_IO_089 */
    mb1_BA3_IO_090_mb1_BC3_IO_080,  /* BA3_IO_090 */
    mb1_BA3_IO_091_mb1_BC3_IO_081,  /* BA3_IO_091 */
    mb1_BA3_IO_092_mb1_BC3_IO_078,  /* BA3_IO_092 */
    mb1_BA3_IO_093_mb1_BC3_IO_079,  /* BA3_IO_093 */
    mb1_BA3_IO_094_mb1_BC3_IO_096,  /* BA3_IO_094 */
    mb1_BA3_IO_095_mb1_BC3_IO_097,  /* BA3_IO_095 */
    mb1_BA3_IO_096_mb1_BC3_IO_094,  /* BA3_IO_096 */
    mb1_BA3_IO_097_mb1_BC3_IO_095,  /* BA3_IO_097 */
    mb1_BA3_IO_098_mb1_BC3_IO_112,  /* BA3_IO_098 */
    mb1_BA3_IO_099_mb1_BC3_IO_113,  /* BA3_IO_099 */
    mb1_BA3_IO_100_mb1_BC3_IO_110,  /* BA3_IO_100 */
    mb1_BA3_IO_101_mb1_BC3_IO_111,  /* BA3_IO_101 */
    mb1_BA3_IO_102_mb1_BC3_IO_088,  /* BA3_IO_102 */
    mb1_BA3_IO_103_mb1_BC3_IO_089,  /* BA3_IO_103 */
    mb1_BA3_IO_104_mb1_BC3_IO_106,  /* BA3_IO_104 */
    mb1_BA3_IO_105_mb1_BC3_IO_107,  /* BA3_IO_105 */

    mb1_BD1_CLKIO_N_0_mb1_BD3_CLKIO_N_7,  /* BD1_CLKIO_N_0 */
    mb1_BD1_CLKIO_N_1_mb1_BD3_CLKIO_N_6,  /* BD1_CLKIO_N_1 */
    mb1_BD1_CLKIO_N_2_mb1_BD3_CLKIO_N_4,  /* BD1_CLKIO_N_2 */
    mb1_BD1_CLKIO_N_3_mb1_BD3_CLKIO_N_3,  /* BD1_CLKIO_N_3 */
    mb1_BD1_CLKIO_N_4_mb1_BD3_CLKIO_N_2,  /* BD1_CLKIO_N_4 */
    mb1_BD1_CLKIO_N_5_mb1_BD3_IO_010,  /* BD1_CLKIO_N_5 */
    mb1_BD1_CLKIO_N_6_mb1_BD3_CLKIO_N_1,  /* BD1_CLKIO_N_6 */
    mb1_BD1_CLKIO_N_7_mb1_BD3_CLKIO_N_0,  /* BD1_CLKIO_N_7 */
    mb1_BD1_CLKIO_P_0_mb1_BD3_CLKIO_P_7,  /* BD1_CLKIO_P_0 */
    mb1_BD1_CLKIO_P_1_mb1_BD3_CLKIO_P_6,  /* BD1_CLKIO_P_1 */
    mb1_BD1_CLKIO_P_2_mb1_BD3_CLKIO_P_4,  /* BD1_CLKIO_P_2 */
    mb1_BD1_CLKIO_P_3_mb1_BD3_CLKIO_P_3,  /* BD1_CLKIO_P_3 */
    mb1_BD1_CLKIO_P_4_mb1_BD3_CLKIO_P_2,  /* BD1_CLKIO_P_4 */
    mb1_BD1_CLKIO_P_5_mb1_BD3_IO_011,  /* BD1_CLKIO_P_5 */
    mb1_BD1_CLKIO_P_6_mb1_BD3_CLKIO_P_1,  /* BD1_CLKIO_P_6 */
    mb1_BD1_CLKIO_P_7_mb1_BD3_CLKIO_P_0,  /* BD1_CLKIO_P_7 */
    mb1_BD1_IO_004_mb1_BD3_IO_006,  /* BD1_IO_004 */
    mb1_BD1_IO_005_mb1_BD3_IO_007,  /* BD1_IO_005 */
    mb1_BD1_IO_006_mb1_BD3_IO_004,  /* BD1_IO_006 */
    mb1_BD1_IO_007_mb1_BD3_IO_005,  /* BD1_IO_007 */
    mb1_BD1_IO_008_mb1_BD3_IO_022,  /* BD1_IO_008 */
    mb1_BD1_IO_009_mb1_BD3_IO_023,  /* BD1_IO_009 */
    mb1_BD1_IO_010_mb1_BD3_CLKIO_N_5,  /* BD1_IO_010 */
    mb1_BD1_IO_011_mb1_BD3_CLKIO_P_5,  /* BD1_IO_011 */
    mb1_BD1_IO_012_mb1_BD3_IO_012,  /* BD1_IO_012 */
    mb1_BD1_IO_013_mb1_BD3_IO_013,  /* BD1_IO_013 */
    mb1_BD1_IO_014_mb1_BD3_IO_016,  /* BD1_IO_014 */
    mb1_BD1_IO_015_mb1_BD3_IO_017,  /* BD1_IO_015 */
    mb1_BD1_IO_016_mb1_BD3_IO_014,  /* BD1_IO_016 */
    mb1_BD1_IO_017_mb1_BD3_IO_015,  /* BD1_IO_017 */
    mb1_BD1_IO_018_mb1_BD3_IO_032,  /* BD1_IO_018 */
    mb1_BD1_IO_019_mb1_BD3_IO_033,  /* BD1_IO_019 */
    mb1_BD1_IO_020_mb1_BD3_IO_030,  /* BD1_IO_020 */
    mb1_BD1_IO_021_mb1_BD3_IO_031,  /* BD1_IO_021 */
    mb1_BD1_IO_022_mb1_BD3_IO_008,  /* BD1_IO_022 */
    mb1_BD1_IO_023_mb1_BD3_IO_009,  /* BD1_IO_023 */
    mb1_BD1_IO_024_mb1_BD3_IO_026,  /* BD1_IO_024 */
    mb1_BD1_IO_025_mb1_BD3_IO_027,  /* BD1_IO_025 */
    mb1_BD1_IO_026_mb1_BD3_IO_024,  /* BD1_IO_026 */
    mb1_BD1_IO_027_mb1_BD3_IO_025,  /* BD1_IO_027 */
    mb1_BD1_IO_028_mb1_BD3_IO_042,  /* BD1_IO_028 */
    mb1_BD1_IO_029_mb1_BD3_IO_043,  /* BD1_IO_029 */
    mb1_BD1_IO_030_mb1_BD3_IO_020,  /* BD1_IO_030 */
    mb1_BD1_IO_031_mb1_BD3_IO_021,  /* BD1_IO_031 */
    mb1_BD1_IO_032_mb1_BD3_IO_018,  /* BD1_IO_032 */
    mb1_BD1_IO_033_mb1_BD3_IO_019,  /* BD1_IO_033 */
    mb1_BD1_IO_034_mb1_BD3_IO_036,  /* BD1_IO_034 */
    mb1_BD1_IO_035_mb1_BD3_IO_037,  /* BD1_IO_035 */
    mb1_BD1_IO_036_mb1_BD3_IO_034,  /* BD1_IO_036 */
    mb1_BD1_IO_037_mb1_BD3_IO_035,  /* BD1_IO_037 */
    mb1_BD1_IO_038_mb1_BD3_IO_052,  /* BD1_IO_038 */
    mb1_BD1_IO_039_mb1_BD3_IO_053,  /* BD1_IO_039 */
    mb1_BD1_IO_040_mb1_BD3_IO_050,  /* BD1_IO_040 */
    mb1_BD1_IO_041_mb1_BD3_IO_051,  /* BD1_IO_041 */
    mb1_BD1_IO_042_mb1_BD3_IO_028,  /* BD1_IO_042 */
    mb1_BD1_IO_043_mb1_BD3_IO_029,  /* BD1_IO_043 */
    mb1_BD1_IO_044_mb1_BD3_IO_046,  /* BD1_IO_044 */
    mb1_BD1_IO_045_mb1_BD3_IO_047,  /* BD1_IO_045 */
    mb1_BD1_IO_046_mb1_BD3_IO_044,  /* BD1_IO_046 */
    mb1_BD1_IO_047_mb1_BD3_IO_045,  /* BD1_IO_047 */
    mb1_BD1_IO_048_mb1_BD3_IO_062,  /* BD1_IO_048 */
    mb1_BD1_IO_049_mb1_BD3_IO_063,  /* BD1_IO_049 */
    mb1_BD1_IO_050_mb1_BD3_IO_040,  /* BD1_IO_050 */
    mb1_BD1_IO_051_mb1_BD3_IO_041,  /* BD1_IO_051 */
    mb1_BD1_IO_052_mb1_BD3_IO_038,  /* BD1_IO_052 */
    mb1_BD1_IO_053_mb1_BD3_IO_039,  /* BD1_IO_053 */
    mb1_BD1_IO_054_mb1_BD3_IO_056,  /* BD1_IO_054 */
    mb1_BD1_IO_055_mb1_BD3_IO_057,  /* BD1_IO_055 */
    mb1_BD1_IO_056_mb1_BD3_IO_054,  /* BD1_IO_056 */
    mb1_BD1_IO_057_mb1_BD3_IO_055,  /* BD1_IO_057 */
    mb1_BD1_IO_058_mb1_BD3_IO_072,  /* BD1_IO_058 */
    mb1_BD1_IO_059_mb1_BD3_IO_073,  /* BD1_IO_059 */
    mb1_BD1_IO_060_mb1_BD3_IO_070,  /* BD1_IO_060 */
    mb1_BD1_IO_061_mb1_BD3_IO_071,  /* BD1_IO_061 */
    mb1_BD1_IO_062_mb1_BD3_IO_048,  /* BD1_IO_062 */
    mb1_BD1_IO_063_mb1_BD3_IO_049,  /* BD1_IO_063 */
    mb1_BD1_IO_064_mb1_BD3_IO_066,  /* BD1_IO_064 */
    mb1_BD1_IO_065_mb1_BD3_IO_067,  /* BD1_IO_065 */
    mb1_BD1_IO_066_mb1_BD3_IO_064,  /* BD1_IO_066 */
    mb1_BD1_IO_067_mb1_BD3_IO_065,  /* BD1_IO_067 */
    mb1_BD1_IO_068_mb1_BD3_IO_082,  /* BD1_IO_068 */
    mb1_BD1_IO_069_mb1_BD3_IO_083,  /* BD1_IO_069 */
    mb1_BD1_IO_070_mb1_BD3_IO_060,  /* BD1_IO_070 */
    mb1_BD1_IO_071_mb1_BD3_IO_061,  /* BD1_IO_071 */
    mb1_BD1_IO_072_mb1_BD3_IO_058,  /* BD1_IO_072 */
    mb1_BD1_IO_073_mb1_BD3_IO_059,  /* BD1_IO_073 */
    mb1_BD1_IO_074_mb1_BD3_IO_076,  /* BD1_IO_074 */
    mb1_BD1_IO_075_mb1_BD3_IO_077,  /* BD1_IO_075 */
    mb1_BD1_IO_076_mb1_BD3_IO_074,  /* BD1_IO_076 */
    mb1_BD1_IO_077_mb1_BD3_IO_075,  /* BD1_IO_077 */
    mb1_BD1_IO_078_mb1_BD3_IO_092,  /* BD1_IO_078 */
    mb1_BD1_IO_079_mb1_BD3_IO_093,  /* BD1_IO_079 */
    mb1_BD1_IO_080_mb1_BD3_IO_090,  /* BD1_IO_080 */
    mb1_BD1_IO_081_mb1_BD3_IO_091,  /* BD1_IO_081 */
    mb1_BD1_IO_082_mb1_BD3_IO_068,  /* BD1_IO_082 */
    mb1_BD1_IO_083_mb1_BD3_IO_069,  /* BD1_IO_083 */
    mb1_BD1_IO_084_mb1_BD3_IO_086,  /* BD1_IO_084 */
    mb1_BD1_IO_085_mb1_BD3_IO_087,  /* BD1_IO_085 */
    mb1_BD1_IO_086_mb1_BD3_IO_084,  /* BD1_IO_086 */
    mb1_BD1_IO_087_mb1_BD3_IO_085,  /* BD1_IO_087 */
    mb1_BD1_IO_088_mb1_BD3_IO_102,  /* BD1_IO_088 */
    mb1_BD1_IO_089_mb1_BD3_IO_103,  /* BD1_IO_089 */
    mb1_BD1_IO_090_mb1_BD3_IO_080,  /* BD1_IO_090 */
    mb1_BD1_IO_091_mb1_BD3_IO_081,  /* BD1_IO_091 */
    mb1_BD1_IO_092_mb1_BD3_IO_078,  /* BD1_IO_092 */
    mb1_BD1_IO_093_mb1_BD3_IO_079,  /* BD1_IO_093 */
    mb1_BD1_IO_094_mb1_BD3_IO_096,  /* BD1_IO_094 */
    mb1_BD1_IO_095_mb1_BD3_IO_097,  /* BD1_IO_095 */
    mb1_BD1_IO_096_mb1_BD3_IO_094,  /* BD1_IO_096 */
    mb1_BD1_IO_097_mb1_BD3_IO_095,  /* BD1_IO_097 */
    mb1_BD1_IO_098_mb1_BD3_IO_112,  /* BD1_IO_098 */
    mb1_BD1_IO_099_mb1_BD3_IO_113,  /* BD1_IO_099 */
    mb1_BD1_IO_100_mb1_BD3_IO_110,  /* BD1_IO_100 */
    mb1_BD1_IO_101_mb1_BD3_IO_111,  /* BD1_IO_101 */
    mb1_BD1_IO_102_mb1_BD3_IO_088,  /* BD1_IO_102 */
    mb1_BD1_IO_103_mb1_BD3_IO_089,  /* BD1_IO_103 */
    mb1_BD1_IO_104_mb1_BD3_IO_106,  /* BD1_IO_104 */
    mb1_BD1_IO_105_mb1_BD3_IO_107
    );

    /* pins which are not connected to an x-board */
    parameter ADDR_W  = 22;
    parameter DQ_PINS = 18;
    parameter GROUPS  = 2;

    output logic               sram0_k_p;
    output logic               sram0_k_n;
    output logic [ADDR_W-1:0]  sram0_a;
    inout  tri   [DQ_PINS-1:0] sram0_dq;
    output logic [GROUPS-1:0]  sram0_bws_n;
    output logic               sram0_rnw;
    output logic               sram0_ld_n;
    output logic               sram0_doff_n;

    output logic               sram1_k_p;
    output logic               sram1_k_n;
    output logic [ADDR_W-1:0]  sram1_a;
    inout  tri   [DQ_PINS-1:0] sram1_dq;
    output logic [GROUPS-1:0]  sram1_bws_n;
    output logic               sram1_rnw;
    output logic               sram1_ld_n;
    output logic               sram1_doff_n;

    output logic               sram2_k_p;
    output logic               sram2_k_n;
    output logic [ADDR_W-1:0]  sram2_a;
    inout  tri   [DQ_PINS-1:0] sram2_dq;
    output logic [GROUPS-1:0]  sram2_bws_n;
    output logic               sram2_rnw;
    output logic               sram2_ld_n;
    output logic               sram2_doff_n;

    output logic               sram3_k_p;
    output logic               sram3_k_n;
    output logic [ADDR_W-1:0]  sram3_a;
    inout  tri   [DQ_PINS-1:0] sram3_dq;
    output logic [GROUPS-1:0]  sram3_bws_n;
    output logic               sram3_rnw;
    output logic               sram3_ld_n;
    output logic               sram3_doff_n;

    `ifdef EN_DDR
        inout wire  [63:0] ddr3_dq;
        inout wire  [7:0]  ddr3_dqs_n;
        inout wire  [7:0]  ddr3_dqs_p;
        output wire [14:0] ddr3_addr;
        output wire [2:0]  ddr3_ba;
        output wire        ddr3_ras_n;
        output wire        ddr3_cas_n;
        output wire        ddr3_we_n;
        output wire        ddr3_reset_n;
        output wire        ddr3_ck_p;
        output wire        ddr3_ck_n;
        output wire        ddr3_cke;
        output wire        ddr3_cs_n;
        output wire [7:0]  ddr3_dm;
        output wire        ddr3_odt;
    `endif

    `ifdef EN_ETH
        input  logic       eth_clk_to_mac;
        input  logic       eth_col_clk_mac_freq;
        input  logic       eth_crs_rgmii_sel0;
        output logic       eth_gtx_clk_tck;
        output logic       eth_mdc;
        inout  tri         eth_mdio;
        input  logic       eth_ninterrupt;
        output logic       eth_nreset;
        input  logic       eth_rx_clk;
        input  logic       eth_rx_dv_rck;
        input  logic       eth_rx_er_rxdv_er;
        input  logic [7:0] eth_rxd;
        input  logic       eth_tx_clk_rgmii_sel1;
        output logic       eth_tx_en_txen_er;
        output logic       eth_tx_er;
        output logic [7:0] eth_txd;
    `endif

    output logic [19:0] dmbi_f2h;
    input  logic [19:0] dmbi_h2f;

    input logic clk0_p;
    input logic clk0_n;
    input logic sync0_p;
    input logic sync0_n;

    input logic clk1_p;
    input logic clk1_n;
    input logic sync1_p;
    input logic sync1_n;

    output logic led_red;
    output logic led_green;
    output logic led_blue;
    output logic led_yellow;

    `ifdef EN_DDR
        input logic clk2_n;
        input logic clk2_p;
    `endif

    /* pins which are connected to motherboard connector BA3 */
    /* and connector BA2 on x-board IC-PDS-CABLE-R1 */
    output wire mb1_BA3_CLKIO_N_0_mb1_BC3_CLKIO_N_7;
    output wire mb1_BA3_CLKIO_N_1_mb1_BC3_CLKIO_N_6;
    output wire mb1_BA3_CLKIO_N_2_mb1_BC3_CLKIO_N_4;
    output wire mb1_BA3_CLKIO_N_3_mb1_BC3_CLKIO_N_3;
    output wire mb1_BA3_CLKIO_N_4_mb1_BC3_CLKIO_N_2;
    output wire mb1_BA3_CLKIO_N_5_mb1_BC3_IO_010;
    output wire mb1_BA3_CLKIO_N_6_mb1_BC3_CLKIO_N_1;
    output wire mb1_BA3_CLKIO_N_7_mb1_BC3_CLKIO_N_0;
    output wire mb1_BA3_CLKIO_P_0_mb1_BC3_CLKIO_P_7;
    output wire mb1_BA3_CLKIO_P_1_mb1_BC3_CLKIO_P_6;
    output wire mb1_BA3_CLKIO_P_2_mb1_BC3_CLKIO_P_4;
    output wire mb1_BA3_CLKIO_P_3_mb1_BC3_CLKIO_P_3;
    output wire mb1_BA3_CLKIO_P_4_mb1_BC3_CLKIO_P_2;
    output wire mb1_BA3_CLKIO_P_5_mb1_BC3_IO_011;
    output wire mb1_BA3_CLKIO_P_6_mb1_BC3_CLKIO_P_1;
    output wire mb1_BA3_CLKIO_P_7_mb1_BC3_CLKIO_P_0;
    output wire mb1_BA3_IO_004_mb1_BC3_IO_006;
    output wire mb1_BA3_IO_005_mb1_BC3_IO_007;
    output wire mb1_BA3_IO_006_mb1_BC3_IO_004;
    output wire mb1_BA3_IO_007_mb1_BC3_IO_005;
    output wire mb1_BA3_IO_008_mb1_BC3_IO_022;
    output wire mb1_BA3_IO_009_mb1_BC3_IO_023;
    output wire mb1_BA3_IO_010_mb1_BC3_CLKIO_N_5;
    output wire mb1_BA3_IO_011_mb1_BC3_CLKIO_P_5;
    output wire mb1_BA3_IO_012_mb1_BC3_IO_012;
    output wire mb1_BA3_IO_013_mb1_BC3_IO_013;
    output wire mb1_BA3_IO_014_mb1_BC3_IO_016;
    output wire mb1_BA3_IO_015_mb1_BC3_IO_017;
    output wire mb1_BA3_IO_016_mb1_BC3_IO_014;
    output wire mb1_BA3_IO_017_mb1_BC3_IO_015;
    output wire mb1_BA3_IO_018_mb1_BC3_IO_032;
    output wire mb1_BA3_IO_019_mb1_BC3_IO_033;
    output wire mb1_BA3_IO_020_mb1_BC3_IO_030;
    output wire mb1_BA3_IO_021_mb1_BC3_IO_031;
    output wire mb1_BA3_IO_022_mb1_BC3_IO_008;
    output wire mb1_BA3_IO_023_mb1_BC3_IO_009;
    output wire mb1_BA3_IO_024_mb1_BC3_IO_026;
    output wire mb1_BA3_IO_025_mb1_BC3_IO_027;
    output wire mb1_BA3_IO_026_mb1_BC3_IO_024;
    output wire mb1_BA3_IO_027_mb1_BC3_IO_025;
    output wire mb1_BA3_IO_028_mb1_BC3_IO_042;
    output wire mb1_BA3_IO_029_mb1_BC3_IO_043;
    output wire mb1_BA3_IO_030_mb1_BC3_IO_020;
    output wire mb1_BA3_IO_031_mb1_BC3_IO_021;
    output wire mb1_BA3_IO_032_mb1_BC3_IO_018;
    output wire mb1_BA3_IO_033_mb1_BC3_IO_019;
    output wire mb1_BA3_IO_034_mb1_BC3_IO_036;
    output wire mb1_BA3_IO_035_mb1_BC3_IO_037;
    output wire mb1_BA3_IO_036_mb1_BC3_IO_034;
    output wire mb1_BA3_IO_037_mb1_BC3_IO_035;
    output wire mb1_BA3_IO_038_mb1_BC3_IO_052;
    output wire mb1_BA3_IO_039_mb1_BC3_IO_053;
    output wire mb1_BA3_IO_040_mb1_BC3_IO_050;
    output wire mb1_BA3_IO_041_mb1_BC3_IO_051;
    output wire mb1_BA3_IO_042_mb1_BC3_IO_028;
    output wire mb1_BA3_IO_043_mb1_BC3_IO_029;
    output wire mb1_BA3_IO_044_mb1_BC3_IO_046;
    output wire mb1_BA3_IO_045_mb1_BC3_IO_047;
    output wire mb1_BA3_IO_046_mb1_BC3_IO_044;

    input wire mb1_BA3_IO_047_mb1_BC3_IO_045;
    input wire mb1_BA3_IO_048_mb1_BC3_IO_062;
    input wire mb1_BA3_IO_049_mb1_BC3_IO_063;
    input wire mb1_BA3_IO_050_mb1_BC3_IO_040;
    input wire mb1_BA3_IO_051_mb1_BC3_IO_041;
    input wire mb1_BA3_IO_052_mb1_BC3_IO_038;
    input wire mb1_BA3_IO_053_mb1_BC3_IO_039;
    input wire mb1_BA3_IO_054_mb1_BC3_IO_056;
    input wire mb1_BA3_IO_055_mb1_BC3_IO_057;
    input wire mb1_BA3_IO_056_mb1_BC3_IO_054;
    input wire mb1_BA3_IO_057_mb1_BC3_IO_055;
    input wire mb1_BA3_IO_058_mb1_BC3_IO_072;
    input wire mb1_BA3_IO_059_mb1_BC3_IO_073;
    input wire mb1_BA3_IO_060_mb1_BC3_IO_070;
    input wire mb1_BA3_IO_061_mb1_BC3_IO_071;
    input wire mb1_BA3_IO_062_mb1_BC3_IO_048;
    input wire mb1_BA3_IO_063_mb1_BC3_IO_049;
    input wire mb1_BA3_IO_064_mb1_BC3_IO_066;
    input wire mb1_BA3_IO_065_mb1_BC3_IO_067;
    input wire mb1_BA3_IO_066_mb1_BC3_IO_064;
    input wire mb1_BA3_IO_067_mb1_BC3_IO_065;
    input wire mb1_BA3_IO_068_mb1_BC3_IO_082;
    input wire mb1_BA3_IO_069_mb1_BC3_IO_083;
    input wire mb1_BA3_IO_070_mb1_BC3_IO_060;
    input wire mb1_BA3_IO_071_mb1_BC3_IO_061;
    input wire mb1_BA3_IO_072_mb1_BC3_IO_058;
    input wire mb1_BA3_IO_073_mb1_BC3_IO_059;
    input wire mb1_BA3_IO_074_mb1_BC3_IO_076;
    input wire mb1_BA3_IO_075_mb1_BC3_IO_077;
    input wire mb1_BA3_IO_076_mb1_BC3_IO_074;
    input wire mb1_BA3_IO_077_mb1_BC3_IO_075;
    input wire mb1_BA3_IO_078_mb1_BC3_IO_092;
    input wire mb1_BA3_IO_079_mb1_BC3_IO_093;
    input wire mb1_BA3_IO_080_mb1_BC3_IO_090;
    input wire mb1_BA3_IO_081_mb1_BC3_IO_091;
    input wire mb1_BA3_IO_082_mb1_BC3_IO_068;
    input wire mb1_BA3_IO_083_mb1_BC3_IO_069;
    input wire mb1_BA3_IO_084_mb1_BC3_IO_086;
    input wire mb1_BA3_IO_085_mb1_BC3_IO_087;
    input wire mb1_BA3_IO_086_mb1_BC3_IO_084;
    input wire mb1_BA3_IO_087_mb1_BC3_IO_085;
    input wire mb1_BA3_IO_088_mb1_BC3_IO_102;
    input wire mb1_BA3_IO_089_mb1_BC3_IO_103;
    input wire mb1_BA3_IO_090_mb1_BC3_IO_080;
    input wire mb1_BA3_IO_091_mb1_BC3_IO_081;
    input wire mb1_BA3_IO_092_mb1_BC3_IO_078;
    input wire mb1_BA3_IO_093_mb1_BC3_IO_079;
    input wire mb1_BA3_IO_094_mb1_BC3_IO_096;
    input wire mb1_BA3_IO_095_mb1_BC3_IO_097;
    input wire mb1_BA3_IO_096_mb1_BC3_IO_094;
    input wire mb1_BA3_IO_097_mb1_BC3_IO_095;
    input wire mb1_BA3_IO_098_mb1_BC3_IO_112;
    input wire mb1_BA3_IO_099_mb1_BC3_IO_113;
    input wire mb1_BA3_IO_100_mb1_BC3_IO_110;
    input wire mb1_BA3_IO_101_mb1_BC3_IO_111;
    input wire mb1_BA3_IO_102_mb1_BC3_IO_088;
    input wire mb1_BA3_IO_103_mb1_BC3_IO_089;
    input wire mb1_BA3_IO_104_mb1_BC3_IO_106;
    input wire mb1_BA3_IO_105_mb1_BC3_IO_107;

    /* pins which are connected to motherboard connector BD1 */
    /* and connector BA2 on x-board IC-PDS-CABLE-R1 */
    output wire mb1_BD1_CLKIO_N_0_mb1_BD3_CLKIO_N_7;
    output wire mb1_BD1_CLKIO_N_1_mb1_BD3_CLKIO_N_6;
    output wire mb1_BD1_CLKIO_N_2_mb1_BD3_CLKIO_N_4;
    output wire mb1_BD1_CLKIO_N_3_mb1_BD3_CLKIO_N_3;
    output wire mb1_BD1_CLKIO_N_4_mb1_BD3_CLKIO_N_2;
    output wire mb1_BD1_CLKIO_N_5_mb1_BD3_IO_010;
    output wire mb1_BD1_CLKIO_N_6_mb1_BD3_CLKIO_N_1;
    output wire mb1_BD1_CLKIO_N_7_mb1_BD3_CLKIO_N_0;
    output wire mb1_BD1_CLKIO_P_0_mb1_BD3_CLKIO_P_7;
    output wire mb1_BD1_CLKIO_P_1_mb1_BD3_CLKIO_P_6;
    output wire mb1_BD1_CLKIO_P_2_mb1_BD3_CLKIO_P_4;
    output wire mb1_BD1_CLKIO_P_3_mb1_BD3_CLKIO_P_3;
    output wire mb1_BD1_CLKIO_P_4_mb1_BD3_CLKIO_P_2;
    output wire mb1_BD1_CLKIO_P_5_mb1_BD3_IO_011;
    output wire mb1_BD1_CLKIO_P_6_mb1_BD3_CLKIO_P_1;
    output wire mb1_BD1_CLKIO_P_7_mb1_BD3_CLKIO_P_0;
    output wire mb1_BD1_IO_004_mb1_BD3_IO_006;
    output wire mb1_BD1_IO_005_mb1_BD3_IO_007;
    output wire mb1_BD1_IO_006_mb1_BD3_IO_004;
    output wire mb1_BD1_IO_007_mb1_BD3_IO_005;
    output wire mb1_BD1_IO_008_mb1_BD3_IO_022;
    output wire mb1_BD1_IO_009_mb1_BD3_IO_023;
    output wire mb1_BD1_IO_010_mb1_BD3_CLKIO_N_5;
    output wire mb1_BD1_IO_011_mb1_BD3_CLKIO_P_5;
    output wire mb1_BD1_IO_012_mb1_BD3_IO_012;
    output wire mb1_BD1_IO_013_mb1_BD3_IO_013;
    output wire mb1_BD1_IO_014_mb1_BD3_IO_016;
    output wire mb1_BD1_IO_015_mb1_BD3_IO_017;
    output wire mb1_BD1_IO_016_mb1_BD3_IO_014;
    output wire mb1_BD1_IO_017_mb1_BD3_IO_015;
    output wire mb1_BD1_IO_018_mb1_BD3_IO_032;
    output wire mb1_BD1_IO_019_mb1_BD3_IO_033;
    output wire mb1_BD1_IO_020_mb1_BD3_IO_030;
    output wire mb1_BD1_IO_021_mb1_BD3_IO_031;
    output wire mb1_BD1_IO_022_mb1_BD3_IO_008;
    output wire mb1_BD1_IO_023_mb1_BD3_IO_009;
    output wire mb1_BD1_IO_024_mb1_BD3_IO_026;
    output wire mb1_BD1_IO_025_mb1_BD3_IO_027;
    output wire mb1_BD1_IO_026_mb1_BD3_IO_024;
    output wire mb1_BD1_IO_027_mb1_BD3_IO_025;
    output wire mb1_BD1_IO_028_mb1_BD3_IO_042;
    output wire mb1_BD1_IO_029_mb1_BD3_IO_043;
    output wire mb1_BD1_IO_030_mb1_BD3_IO_020;
    output wire mb1_BD1_IO_031_mb1_BD3_IO_021;
    output wire mb1_BD1_IO_032_mb1_BD3_IO_018;
    output wire mb1_BD1_IO_033_mb1_BD3_IO_019;
    output wire mb1_BD1_IO_034_mb1_BD3_IO_036;
    output wire mb1_BD1_IO_035_mb1_BD3_IO_037;
    output wire mb1_BD1_IO_036_mb1_BD3_IO_034;
    output wire mb1_BD1_IO_037_mb1_BD3_IO_035;
    output wire mb1_BD1_IO_038_mb1_BD3_IO_052;
    output wire mb1_BD1_IO_039_mb1_BD3_IO_053;
    output wire mb1_BD1_IO_040_mb1_BD3_IO_050;
    output wire mb1_BD1_IO_041_mb1_BD3_IO_051;
    output wire mb1_BD1_IO_042_mb1_BD3_IO_028;
    output wire mb1_BD1_IO_043_mb1_BD3_IO_029;
    output wire mb1_BD1_IO_044_mb1_BD3_IO_046;
    output wire mb1_BD1_IO_045_mb1_BD3_IO_047;
    output wire mb1_BD1_IO_046_mb1_BD3_IO_044;

    input wire mb1_BD1_IO_047_mb1_BD3_IO_045;
    input wire mb1_BD1_IO_048_mb1_BD3_IO_062;
    input wire mb1_BD1_IO_049_mb1_BD3_IO_063;
    input wire mb1_BD1_IO_050_mb1_BD3_IO_040;
    input wire mb1_BD1_IO_051_mb1_BD3_IO_041;
    input wire mb1_BD1_IO_052_mb1_BD3_IO_038;
    input wire mb1_BD1_IO_053_mb1_BD3_IO_039;
    input wire mb1_BD1_IO_054_mb1_BD3_IO_056;
    input wire mb1_BD1_IO_055_mb1_BD3_IO_057;
    input wire mb1_BD1_IO_056_mb1_BD3_IO_054;
    input wire mb1_BD1_IO_057_mb1_BD3_IO_055;
    input wire mb1_BD1_IO_058_mb1_BD3_IO_072;
    input wire mb1_BD1_IO_059_mb1_BD3_IO_073;
    input wire mb1_BD1_IO_060_mb1_BD3_IO_070;
    input wire mb1_BD1_IO_061_mb1_BD3_IO_071;
    input wire mb1_BD1_IO_062_mb1_BD3_IO_048;
    input wire mb1_BD1_IO_063_mb1_BD3_IO_049;
    input wire mb1_BD1_IO_064_mb1_BD3_IO_066;
    input wire mb1_BD1_IO_065_mb1_BD3_IO_067;
    input wire mb1_BD1_IO_066_mb1_BD3_IO_064;
    input wire mb1_BD1_IO_067_mb1_BD3_IO_065;
    input wire mb1_BD1_IO_068_mb1_BD3_IO_082;
    input wire mb1_BD1_IO_069_mb1_BD3_IO_083;
    input wire mb1_BD1_IO_070_mb1_BD3_IO_060;
    input wire mb1_BD1_IO_071_mb1_BD3_IO_061;
    input wire mb1_BD1_IO_072_mb1_BD3_IO_058;
    input wire mb1_BD1_IO_073_mb1_BD3_IO_059;
    input wire mb1_BD1_IO_074_mb1_BD3_IO_076;
    input wire mb1_BD1_IO_075_mb1_BD3_IO_077;
    input wire mb1_BD1_IO_076_mb1_BD3_IO_074;
    input wire mb1_BD1_IO_077_mb1_BD3_IO_075;
    input wire mb1_BD1_IO_078_mb1_BD3_IO_092;
    input wire mb1_BD1_IO_079_mb1_BD3_IO_093;
    input wire mb1_BD1_IO_080_mb1_BD3_IO_090;
    input wire mb1_BD1_IO_081_mb1_BD3_IO_091;
    input wire mb1_BD1_IO_082_mb1_BD3_IO_068;
    input wire mb1_BD1_IO_083_mb1_BD3_IO_069;
    input wire mb1_BD1_IO_084_mb1_BD3_IO_086;
    input wire mb1_BD1_IO_085_mb1_BD3_IO_087;
    input wire mb1_BD1_IO_086_mb1_BD3_IO_084;
    input wire mb1_BD1_IO_087_mb1_BD3_IO_085;
    input wire mb1_BD1_IO_088_mb1_BD3_IO_102;
    input wire mb1_BD1_IO_089_mb1_BD3_IO_103;
    input wire mb1_BD1_IO_090_mb1_BD3_IO_080;
    input wire mb1_BD1_IO_091_mb1_BD3_IO_081;
    input wire mb1_BD1_IO_092_mb1_BD3_IO_078;
    input wire mb1_BD1_IO_093_mb1_BD3_IO_079;
    input wire mb1_BD1_IO_094_mb1_BD3_IO_096;
    input wire mb1_BD1_IO_095_mb1_BD3_IO_097;
    input wire mb1_BD1_IO_096_mb1_BD3_IO_094;
    input wire mb1_BD1_IO_097_mb1_BD3_IO_095;
    input wire mb1_BD1_IO_098_mb1_BD3_IO_112;
    input wire mb1_BD1_IO_099_mb1_BD3_IO_113;
    input wire mb1_BD1_IO_100_mb1_BD3_IO_110;
    input wire mb1_BD1_IO_101_mb1_BD3_IO_111;
    input wire mb1_BD1_IO_102_mb1_BD3_IO_088;
    input wire mb1_BD1_IO_103_mb1_BD3_IO_089;
    input wire mb1_BD1_IO_104_mb1_BD3_IO_106;
    input wire mb1_BD1_IO_105_mb1_BD3_IO_107;

    localparam TX_PINS = 59;
    localparam RX_PINS = 59;

    wire [TX_PINS-1:0] tx_pin;
    wire [RX_PINS-1:0] rx_pin;

    assign mb1_BA3_CLKIO_N_0_mb1_BC3_CLKIO_N_7 = tx_pin[0];
    assign mb1_BA3_CLKIO_N_1_mb1_BC3_CLKIO_N_6 = tx_pin[1];
    assign mb1_BA3_CLKIO_N_2_mb1_BC3_CLKIO_N_4 = tx_pin[2];
    assign mb1_BA3_CLKIO_N_3_mb1_BC3_CLKIO_N_3 = tx_pin[3];
    assign mb1_BA3_CLKIO_N_4_mb1_BC3_CLKIO_N_2 = tx_pin[4];
    assign mb1_BA3_CLKIO_N_5_mb1_BC3_IO_010 = tx_pin[5];
    assign mb1_BA3_CLKIO_N_6_mb1_BC3_CLKIO_N_1 = tx_pin[6];
    assign mb1_BA3_CLKIO_N_7_mb1_BC3_CLKIO_N_0 = tx_pin[7];
    assign mb1_BA3_CLKIO_P_0_mb1_BC3_CLKIO_P_7 = tx_pin[8];
    assign mb1_BA3_CLKIO_P_1_mb1_BC3_CLKIO_P_6 = tx_pin[9];
    assign mb1_BA3_CLKIO_P_2_mb1_BC3_CLKIO_P_4 = tx_pin[10];
    assign mb1_BA3_CLKIO_P_3_mb1_BC3_CLKIO_P_3 = tx_pin[11];
    assign mb1_BA3_CLKIO_P_4_mb1_BC3_CLKIO_P_2 = tx_pin[12];
    assign mb1_BA3_CLKIO_P_5_mb1_BC3_IO_011 = tx_pin[13];
    assign mb1_BA3_CLKIO_P_6_mb1_BC3_CLKIO_P_1 = tx_pin[14];
    assign mb1_BA3_CLKIO_P_7_mb1_BC3_CLKIO_P_0 = tx_pin[15];
    assign mb1_BA3_IO_004_mb1_BC3_IO_006 = tx_pin[16];
    assign mb1_BA3_IO_005_mb1_BC3_IO_007 = tx_pin[17];
    assign mb1_BA3_IO_006_mb1_BC3_IO_004 = tx_pin[18];
    assign mb1_BA3_IO_007_mb1_BC3_IO_005 = tx_pin[19];
    assign mb1_BA3_IO_008_mb1_BC3_IO_022 = tx_pin[20];
    assign mb1_BA3_IO_009_mb1_BC3_IO_023 = tx_pin[21];
    assign mb1_BA3_IO_010_mb1_BC3_CLKIO_N_5 = tx_pin[22];
    assign mb1_BA3_IO_011_mb1_BC3_CLKIO_P_5 = tx_pin[23];
    assign mb1_BA3_IO_012_mb1_BC3_IO_012 = tx_pin[24];
    assign mb1_BA3_IO_013_mb1_BC3_IO_013 = tx_pin[25];
    assign mb1_BA3_IO_014_mb1_BC3_IO_016 = tx_pin[26];
    assign mb1_BA3_IO_015_mb1_BC3_IO_017 = tx_pin[27];
    assign mb1_BA3_IO_016_mb1_BC3_IO_014 = tx_pin[28];
    assign mb1_BA3_IO_017_mb1_BC3_IO_015 = tx_pin[29];
    assign mb1_BA3_IO_018_mb1_BC3_IO_032 = tx_pin[30];
    assign mb1_BA3_IO_019_mb1_BC3_IO_033 = tx_pin[31];
    assign mb1_BA3_IO_020_mb1_BC3_IO_030 = tx_pin[32];
    assign mb1_BA3_IO_021_mb1_BC3_IO_031 = tx_pin[33];
    assign mb1_BA3_IO_022_mb1_BC3_IO_008 = tx_pin[34];
    assign mb1_BA3_IO_023_mb1_BC3_IO_009 = tx_pin[35];
    assign mb1_BA3_IO_024_mb1_BC3_IO_026 = tx_pin[36];
    assign mb1_BA3_IO_025_mb1_BC3_IO_027 = tx_pin[37];
    assign mb1_BA3_IO_026_mb1_BC3_IO_024 = tx_pin[38];
    assign mb1_BA3_IO_027_mb1_BC3_IO_025 = tx_pin[39];
    assign mb1_BA3_IO_028_mb1_BC3_IO_042 = tx_pin[40];
    assign mb1_BA3_IO_029_mb1_BC3_IO_043 = tx_pin[41];
    assign mb1_BA3_IO_030_mb1_BC3_IO_020 = tx_pin[42];
    assign mb1_BA3_IO_031_mb1_BC3_IO_021 = tx_pin[43];
    assign mb1_BA3_IO_032_mb1_BC3_IO_018 = tx_pin[44];
    assign mb1_BA3_IO_033_mb1_BC3_IO_019 = tx_pin[45];
    assign mb1_BA3_IO_034_mb1_BC3_IO_036 = tx_pin[46];
    assign mb1_BA3_IO_035_mb1_BC3_IO_037 = tx_pin[47];
    assign mb1_BA3_IO_036_mb1_BC3_IO_034 = tx_pin[48];
    assign mb1_BA3_IO_037_mb1_BC3_IO_035 = tx_pin[49];
    assign mb1_BA3_IO_038_mb1_BC3_IO_052 = tx_pin[50];
    assign mb1_BA3_IO_039_mb1_BC3_IO_053 = tx_pin[51];
    assign mb1_BA3_IO_040_mb1_BC3_IO_050 = tx_pin[52];
    assign mb1_BA3_IO_041_mb1_BC3_IO_051 = tx_pin[53];
    assign mb1_BA3_IO_042_mb1_BC3_IO_028 = tx_pin[54];
    assign mb1_BA3_IO_043_mb1_BC3_IO_029 = tx_pin[55];
    assign mb1_BA3_IO_044_mb1_BC3_IO_046 = tx_pin[56];
    assign mb1_BA3_IO_045_mb1_BC3_IO_047 = tx_pin[57];
    assign mb1_BA3_IO_046_mb1_BC3_IO_044 = tx_pin[58];

    assign rx_pin[0] = mb1_BA3_IO_047_mb1_BC3_IO_045;
    assign rx_pin[1] = mb1_BA3_IO_048_mb1_BC3_IO_062;
    assign rx_pin[2] = mb1_BA3_IO_049_mb1_BC3_IO_063;
    assign rx_pin[3] = mb1_BA3_IO_050_mb1_BC3_IO_040;
    assign rx_pin[4] = mb1_BA3_IO_051_mb1_BC3_IO_041;
    assign rx_pin[5] = mb1_BA3_IO_052_mb1_BC3_IO_038;
    assign rx_pin[6] = mb1_BA3_IO_053_mb1_BC3_IO_039;
    assign rx_pin[7] = mb1_BA3_IO_054_mb1_BC3_IO_056;
    assign rx_pin[8] = mb1_BA3_IO_055_mb1_BC3_IO_057;
    assign rx_pin[9] = mb1_BA3_IO_056_mb1_BC3_IO_054;
    assign rx_pin[10] = mb1_BA3_IO_057_mb1_BC3_IO_055;
    assign rx_pin[11] = mb1_BA3_IO_058_mb1_BC3_IO_072;
    assign rx_pin[12] = mb1_BA3_IO_059_mb1_BC3_IO_073;
    assign rx_pin[13] = mb1_BA3_IO_060_mb1_BC3_IO_070;
    assign rx_pin[14] = mb1_BA3_IO_061_mb1_BC3_IO_071;
    assign rx_pin[15] = mb1_BA3_IO_062_mb1_BC3_IO_048;
    assign rx_pin[16] = mb1_BA3_IO_063_mb1_BC3_IO_049;
    assign rx_pin[17] = mb1_BA3_IO_064_mb1_BC3_IO_066;
    assign rx_pin[18] = mb1_BA3_IO_065_mb1_BC3_IO_067;
    assign rx_pin[19] = mb1_BA3_IO_066_mb1_BC3_IO_064;
    assign rx_pin[20] = mb1_BA3_IO_067_mb1_BC3_IO_065;
    assign rx_pin[21] = mb1_BA3_IO_068_mb1_BC3_IO_082;
    assign rx_pin[22] = mb1_BA3_IO_069_mb1_BC3_IO_083;
    assign rx_pin[23] = mb1_BA3_IO_070_mb1_BC3_IO_060;
    assign rx_pin[24] = mb1_BA3_IO_071_mb1_BC3_IO_061;
    assign rx_pin[25] = mb1_BA3_IO_072_mb1_BC3_IO_058;
    assign rx_pin[26] = mb1_BA3_IO_073_mb1_BC3_IO_059;
    assign rx_pin[27] = mb1_BA3_IO_074_mb1_BC3_IO_076;
    assign rx_pin[28] = mb1_BA3_IO_075_mb1_BC3_IO_077;
    assign rx_pin[29] = mb1_BA3_IO_076_mb1_BC3_IO_074;
    assign rx_pin[30] = mb1_BA3_IO_077_mb1_BC3_IO_075;
    assign rx_pin[31] = mb1_BA3_IO_078_mb1_BC3_IO_092;
    assign rx_pin[32] = mb1_BA3_IO_079_mb1_BC3_IO_093;
    assign rx_pin[33] = mb1_BA3_IO_080_mb1_BC3_IO_090;
    assign rx_pin[34] = mb1_BA3_IO_081_mb1_BC3_IO_091;
    assign rx_pin[35] = mb1_BA3_IO_082_mb1_BC3_IO_068;
    assign rx_pin[36] = mb1_BA3_IO_083_mb1_BC3_IO_069;
    assign rx_pin[37] = mb1_BA3_IO_084_mb1_BC3_IO_086;
    assign rx_pin[38] = mb1_BA3_IO_085_mb1_BC3_IO_087;
    assign rx_pin[39] = mb1_BA3_IO_086_mb1_BC3_IO_084;
    assign rx_pin[40] = mb1_BA3_IO_087_mb1_BC3_IO_085;
    assign rx_pin[41] = mb1_BA3_IO_088_mb1_BC3_IO_102;
    assign rx_pin[42] = mb1_BA3_IO_089_mb1_BC3_IO_103;
    assign rx_pin[43] = mb1_BA3_IO_090_mb1_BC3_IO_080;
    assign rx_pin[44] = mb1_BA3_IO_091_mb1_BC3_IO_081;
    assign rx_pin[45] = mb1_BA3_IO_092_mb1_BC3_IO_078;
    assign rx_pin[46] = mb1_BA3_IO_093_mb1_BC3_IO_079;
    assign rx_pin[47] = mb1_BA3_IO_094_mb1_BC3_IO_096;
    assign rx_pin[48] = mb1_BA3_IO_095_mb1_BC3_IO_097;
    assign rx_pin[49] = mb1_BA3_IO_096_mb1_BC3_IO_094;
    assign rx_pin[50] = mb1_BA3_IO_097_mb1_BC3_IO_095;
    assign rx_pin[51] = mb1_BA3_IO_098_mb1_BC3_IO_112;
    assign rx_pin[52] = mb1_BA3_IO_099_mb1_BC3_IO_113;
    assign rx_pin[53] = mb1_BA3_IO_100_mb1_BC3_IO_110;
    assign rx_pin[54] = mb1_BA3_IO_101_mb1_BC3_IO_111;
    assign rx_pin[55] = mb1_BA3_IO_102_mb1_BC3_IO_088;
    assign rx_pin[56] = mb1_BA3_IO_103_mb1_BC3_IO_089;
    assign rx_pin[57] = mb1_BA3_IO_104_mb1_BC3_IO_106;
    assign rx_pin[58] = mb1_BA3_IO_105_mb1_BC3_IO_107;

    wire [TX_PINS-1:0] tx2_pin;
    wire [RX_PINS-1:0] rx2_pin;

    assign mb1_BD1_CLKIO_N_0_mb1_BD3_CLKIO_N_7 = tx2_pin[0];
    assign mb1_BD1_CLKIO_N_1_mb1_BD3_CLKIO_N_6 = tx2_pin[1];
    assign mb1_BD1_CLKIO_N_2_mb1_BD3_CLKIO_N_4 = tx2_pin[2];
    assign mb1_BD1_CLKIO_N_3_mb1_BD3_CLKIO_N_3 = tx2_pin[3];
    assign mb1_BD1_CLKIO_N_4_mb1_BD3_CLKIO_N_2 = tx2_pin[4];
    assign mb1_BD1_CLKIO_N_5_mb1_BD3_IO_010 = tx2_pin[5];
    assign mb1_BD1_CLKIO_N_6_mb1_BD3_CLKIO_N_1 = tx2_pin[6];
    assign mb1_BD1_CLKIO_N_7_mb1_BD3_CLKIO_N_0 = tx2_pin[7];
    assign mb1_BD1_CLKIO_P_0_mb1_BD3_CLKIO_P_7 = tx2_pin[8];
    assign mb1_BD1_CLKIO_P_1_mb1_BD3_CLKIO_P_6 = tx2_pin[9];
    assign mb1_BD1_CLKIO_P_2_mb1_BD3_CLKIO_P_4 = tx2_pin[10];
    assign mb1_BD1_CLKIO_P_3_mb1_BD3_CLKIO_P_3 = tx2_pin[11];
    assign mb1_BD1_CLKIO_P_4_mb1_BD3_CLKIO_P_2 = tx2_pin[12];
    assign mb1_BD1_CLKIO_P_5_mb1_BD3_IO_011 = tx2_pin[13];
    assign mb1_BD1_CLKIO_P_6_mb1_BD3_CLKIO_P_1 = tx2_pin[14];
    assign mb1_BD1_CLKIO_P_7_mb1_BD3_CLKIO_P_0 = tx2_pin[15];
    assign mb1_BD1_IO_004_mb1_BD3_IO_006 = tx2_pin[16];
    assign mb1_BD1_IO_005_mb1_BD3_IO_007 = tx2_pin[17];
    assign mb1_BD1_IO_006_mb1_BD3_IO_004 = tx2_pin[18];
    assign mb1_BD1_IO_007_mb1_BD3_IO_005 = tx2_pin[19];
    assign mb1_BD1_IO_008_mb1_BD3_IO_022 = tx2_pin[20];
    assign mb1_BD1_IO_009_mb1_BD3_IO_023 = tx2_pin[21];
    assign mb1_BD1_IO_010_mb1_BD3_CLKIO_N_5 = tx2_pin[22];
    assign mb1_BD1_IO_011_mb1_BD3_CLKIO_P_5 = tx2_pin[23];
    assign mb1_BD1_IO_012_mb1_BD3_IO_012 = tx2_pin[24];
    assign mb1_BD1_IO_013_mb1_BD3_IO_013 = tx2_pin[25];
    assign mb1_BD1_IO_014_mb1_BD3_IO_016 = tx2_pin[26];
    assign mb1_BD1_IO_015_mb1_BD3_IO_017 = tx2_pin[27];
    assign mb1_BD1_IO_016_mb1_BD3_IO_014 = tx2_pin[28];
    assign mb1_BD1_IO_017_mb1_BD3_IO_015 = tx2_pin[29];
    assign mb1_BD1_IO_018_mb1_BD3_IO_032 = tx2_pin[30];
    assign mb1_BD1_IO_019_mb1_BD3_IO_033 = tx2_pin[31];
    assign mb1_BD1_IO_020_mb1_BD3_IO_030 = tx2_pin[32];
    assign mb1_BD1_IO_021_mb1_BD3_IO_031 = tx2_pin[33];
    assign mb1_BD1_IO_022_mb1_BD3_IO_008 = tx2_pin[34];
    assign mb1_BD1_IO_023_mb1_BD3_IO_009 = tx2_pin[35];
    assign mb1_BD1_IO_024_mb1_BD3_IO_026 = tx2_pin[36];
    assign mb1_BD1_IO_025_mb1_BD3_IO_027 = tx2_pin[37];
    assign mb1_BD1_IO_026_mb1_BD3_IO_024 = tx2_pin[38];
    assign mb1_BD1_IO_027_mb1_BD3_IO_025 = tx2_pin[39];
    assign mb1_BD1_IO_028_mb1_BD3_IO_042 = tx2_pin[40];
    assign mb1_BD1_IO_029_mb1_BD3_IO_043 = tx2_pin[41];
    assign mb1_BD1_IO_030_mb1_BD3_IO_020 = tx2_pin[42];
    assign mb1_BD1_IO_031_mb1_BD3_IO_021 = tx2_pin[43];
    assign mb1_BD1_IO_032_mb1_BD3_IO_018 = tx2_pin[44];
    assign mb1_BD1_IO_033_mb1_BD3_IO_019 = tx2_pin[45];
    assign mb1_BD1_IO_034_mb1_BD3_IO_036 = tx2_pin[46];
    assign mb1_BD1_IO_035_mb1_BD3_IO_037 = tx2_pin[47];
    assign mb1_BD1_IO_036_mb1_BD3_IO_034 = tx2_pin[48];
    assign mb1_BD1_IO_037_mb1_BD3_IO_035 = tx2_pin[49];
    assign mb1_BD1_IO_038_mb1_BD3_IO_052 = tx2_pin[50];
    assign mb1_BD1_IO_039_mb1_BD3_IO_053 = tx2_pin[51];
    assign mb1_BD1_IO_040_mb1_BD3_IO_050 = tx2_pin[52];
    assign mb1_BD1_IO_041_mb1_BD3_IO_051 = tx2_pin[53];
    assign mb1_BD1_IO_042_mb1_BD3_IO_028 = tx2_pin[54];
    assign mb1_BD1_IO_043_mb1_BD3_IO_029 = tx2_pin[55];
    assign mb1_BD1_IO_044_mb1_BD3_IO_046 = tx2_pin[56];
    assign mb1_BD1_IO_045_mb1_BD3_IO_047 = tx2_pin[57];
    assign mb1_BD1_IO_046_mb1_BD3_IO_044 = tx2_pin[58];

    assign rx2_pin[0] = mb1_BD1_IO_047_mb1_BD3_IO_045;
    assign rx2_pin[1] = mb1_BD1_IO_048_mb1_BD3_IO_062;
    assign rx2_pin[2] = mb1_BD1_IO_049_mb1_BD3_IO_063;
    assign rx2_pin[3] = mb1_BD1_IO_050_mb1_BD3_IO_040;
    assign rx2_pin[4] = mb1_BD1_IO_051_mb1_BD3_IO_041;
    assign rx2_pin[5] = mb1_BD1_IO_052_mb1_BD3_IO_038;
    assign rx2_pin[6] = mb1_BD1_IO_053_mb1_BD3_IO_039;
    assign rx2_pin[7] = mb1_BD1_IO_054_mb1_BD3_IO_056;
    assign rx2_pin[8] = mb1_BD1_IO_055_mb1_BD3_IO_057;
    assign rx2_pin[9] = mb1_BD1_IO_056_mb1_BD3_IO_054;
    assign rx2_pin[10] = mb1_BD1_IO_057_mb1_BD3_IO_055;
    assign rx2_pin[11] = mb1_BD1_IO_058_mb1_BD3_IO_072;
    assign rx2_pin[12] = mb1_BD1_IO_059_mb1_BD3_IO_073;
    assign rx2_pin[13] = mb1_BD1_IO_060_mb1_BD3_IO_070;
    assign rx2_pin[14] = mb1_BD1_IO_061_mb1_BD3_IO_071;
    assign rx2_pin[15] = mb1_BD1_IO_062_mb1_BD3_IO_048;
    assign rx2_pin[16] = mb1_BD1_IO_063_mb1_BD3_IO_049;
    assign rx2_pin[17] = mb1_BD1_IO_064_mb1_BD3_IO_066;
    assign rx2_pin[18] = mb1_BD1_IO_065_mb1_BD3_IO_067;
    assign rx2_pin[19] = mb1_BD1_IO_066_mb1_BD3_IO_064;
    assign rx2_pin[20] = mb1_BD1_IO_067_mb1_BD3_IO_065;
    assign rx2_pin[21] = mb1_BD1_IO_068_mb1_BD3_IO_082;
    assign rx2_pin[22] = mb1_BD1_IO_069_mb1_BD3_IO_083;
    assign rx2_pin[23] = mb1_BD1_IO_070_mb1_BD3_IO_060;
    assign rx2_pin[24] = mb1_BD1_IO_071_mb1_BD3_IO_061;
    assign rx2_pin[25] = mb1_BD1_IO_072_mb1_BD3_IO_058;
    assign rx2_pin[26] = mb1_BD1_IO_073_mb1_BD3_IO_059;
    assign rx2_pin[27] = mb1_BD1_IO_074_mb1_BD3_IO_076;
    assign rx2_pin[28] = mb1_BD1_IO_075_mb1_BD3_IO_077;
    assign rx2_pin[29] = mb1_BD1_IO_076_mb1_BD3_IO_074;
    assign rx2_pin[30] = mb1_BD1_IO_077_mb1_BD3_IO_075;
    assign rx2_pin[31] = mb1_BD1_IO_078_mb1_BD3_IO_092;
    assign rx2_pin[32] = mb1_BD1_IO_079_mb1_BD3_IO_093;
    assign rx2_pin[33] = mb1_BD1_IO_080_mb1_BD3_IO_090;
    assign rx2_pin[34] = mb1_BD1_IO_081_mb1_BD3_IO_091;
    assign rx2_pin[35] = mb1_BD1_IO_082_mb1_BD3_IO_068;
    assign rx2_pin[36] = mb1_BD1_IO_083_mb1_BD3_IO_069;
    assign rx2_pin[37] = mb1_BD1_IO_084_mb1_BD3_IO_086;
    assign rx2_pin[38] = mb1_BD1_IO_085_mb1_BD3_IO_087;
    assign rx2_pin[39] = mb1_BD1_IO_086_mb1_BD3_IO_084;
    assign rx2_pin[40] = mb1_BD1_IO_087_mb1_BD3_IO_085;
    assign rx2_pin[41] = mb1_BD1_IO_088_mb1_BD3_IO_102;
    assign rx2_pin[42] = mb1_BD1_IO_089_mb1_BD3_IO_103;
    assign rx2_pin[43] = mb1_BD1_IO_090_mb1_BD3_IO_080;
    assign rx2_pin[44] = mb1_BD1_IO_091_mb1_BD3_IO_081;
    assign rx2_pin[45] = mb1_BD1_IO_092_mb1_BD3_IO_078;
    assign rx2_pin[46] = mb1_BD1_IO_093_mb1_BD3_IO_079;
    assign rx2_pin[47] = mb1_BD1_IO_094_mb1_BD3_IO_096;
    assign rx2_pin[48] = mb1_BD1_IO_095_mb1_BD3_IO_097;
    assign rx2_pin[49] = mb1_BD1_IO_096_mb1_BD3_IO_094;
    assign rx2_pin[50] = mb1_BD1_IO_097_mb1_BD3_IO_095;
    assign rx2_pin[51] = mb1_BD1_IO_098_mb1_BD3_IO_112;
    assign rx2_pin[52] = mb1_BD1_IO_099_mb1_BD3_IO_113;
    assign rx2_pin[53] = mb1_BD1_IO_100_mb1_BD3_IO_110;
    assign rx2_pin[54] = mb1_BD1_IO_101_mb1_BD3_IO_111;
    assign rx2_pin[55] = mb1_BD1_IO_102_mb1_BD3_IO_088;
    assign rx2_pin[56] = mb1_BD1_IO_103_mb1_BD3_IO_089;
    assign rx2_pin[57] = mb1_BD1_IO_104_mb1_BD3_IO_106;
    assign rx2_pin[58] = mb1_BD1_IO_105_mb1_BD3_IO_107;

    top #(
        .FPGA(TC3),
        .fpga_x(0),
        .fpga_y(1))
    top_inst (
        .clk0_p(clk0_p),
        .clk0_n(clk0_n),

        .sync0_p(sync0_p),
        .sync0_n(sync0_n),

        .dmbi_h2f(dmbi_h2f),
        .dmbi_f2h(dmbi_f2h),

        .tx_pin(tx_pin),
        .rx_pin(rx_pin),

        .tx2_pin(tx2_pin),
        .rx2_pin(rx2_pin),

        .clk1_p(clk1_p),
        .clk1_n(clk1_n),

        .sync1_p(sync1_p),
        .sync1_n(sync1_n),

        .led_red(led_red),
        .led_green(led_green),
        .led_blue(led_blue),
        .led_yellow(led_yellow),

        `ifdef EN_DDR
            .clk2_p(clk2_p),
            .clk2_n(clk2_n),
        `endif

        // SSRAM interface
        .sram0_k_p(sram0_k_p),
        .sram0_k_n(sram0_k_n),
        .sram0_a(sram0_a),
        .sram0_dq(sram0_dq),
        .sram0_bws_n(sram0_bws_n),
        .sram0_rnw(sram0_rnw),
        .sram0_ld_n(sram0_ld_n),
        .sram0_doff_n(sram0_doff_n),

        .sram1_k_p(sram1_k_p),
        .sram1_k_n(sram1_k_n),
        .sram1_a(sram1_a),
        .sram1_dq(sram1_dq),
        .sram1_bws_n(sram1_bws_n),
        .sram1_rnw(sram1_rnw),
        .sram1_ld_n(sram1_ld_n),
        .sram1_doff_n(sram1_doff_n),

        .sram2_k_p(sram2_k_p),
        .sram2_k_n(sram2_k_n),
        .sram2_a(sram2_a),
        .sram2_dq(sram2_dq),
        .sram2_bws_n(sram2_bws_n),
        .sram2_rnw(sram2_rnw),
        .sram2_ld_n(sram2_ld_n),
        .sram2_doff_n(sram2_doff_n),

        .sram3_k_p(sram3_k_p),
        .sram3_k_n(sram3_k_n),
        .sram3_a(sram3_a),
        .sram3_dq(sram3_dq),
        .sram3_bws_n(sram3_bws_n),
        .sram3_rnw(sram3_rnw),
        .sram3_ld_n(sram3_ld_n),
        .sram3_doff_n(sram3_doff_n)

        `ifdef EN_DDR
            ,
            .ddr3_dq(ddr3_dq),
            .ddr3_dqs_p(ddr3_dqs_p),
            .ddr3_dqs_n(ddr3_dqs_n),
            .ddr3_addr(ddr3_addr),
            .ddr3_ba(ddr3_ba),
            .ddr3_ras_n(ddr3_ras_n),
            .ddr3_cas_n(ddr3_cas_n),
            .ddr3_we_n(ddr3_we_n),
            .ddr3_reset_n(ddr3_reset_n),
            .ddr3_ck_p(ddr3_ck_p),
            .ddr3_ck_n(ddr3_ck_n),
            .ddr3_cke(ddr3_cke),
            .ddr3_cs_n(ddr3_cs_n),
            .ddr3_dm(ddr3_dm),
            .ddr3_odt(ddr3_odt)
        `endif

        `ifdef EN_ETH
            ,
            .eth_clk_to_mac(eth_clk_to_mac),
            .eth_col_clk_mac_freq(eth_col_clk_mac_freq),
            .eth_crs_rgmii_sel0(eth_crs_rgmii_sel0),
            .eth_gtx_clk_tck(eth_gtx_clk_tck),
            .eth_mdc(eth_mdc),
            .eth_mdio(eth_mdio),
            .eth_ninterrupt(eth_ninterrupt),
            .eth_nreset(eth_nreset),
            .eth_rx_clk(eth_rx_clk),
            .eth_rx_dv_rck(eth_rx_dv_rck),
            .eth_rx_er_rxdv_er(eth_rx_er_rxdv_er),
            .eth_rxd(eth_rxd),
            .eth_tx_clk_rgmii_sel1(eth_tx_clk_rgmii_sel1),
            .eth_tx_en_txen_er(eth_tx_en_txen_er),
            .eth_tx_er(eth_tx_er),
            .eth_txd(eth_txd)
        `endif
    );
endmodule
