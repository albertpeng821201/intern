/* (c) Copyright 2012-2016 PRO DESIGN Electronic GmbH.                     */
/* All rights reserved.                                                    */
/*                                                                         */
/* This file is owned and controlled by ProDesign and must be used solely  */
/* for design, simulation, implementation and creation of design files     */
/* limited to profpga systems or technologies. Use with non-profpga        */
/* systems or technologies is expressly prohibited and immediately         */
/* terminates your license.                                                */
/*                                                                         */
/* PRODESIGN IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY */
/* FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR PRODESIGN SYSTEMS. BY  */
/* PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             */
/* IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, PRODESIGN IS   */
/* MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      */
/* CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       */
/* RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION. PRODESIGN EXPRESSLY     */
/* DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   */
/* IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          */
/* REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         */
/* INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   */
/* PARTICULAR PURPOSE.                                                     */
/*                                                                         */
/* ProDesign products are not intended for use in life support appliances, */
/* devices, or systems. Use in such applications are expressly             */
/* prohibited.                                                             */
/*                                                                         */
/* This file was generated by profpga_brdgen version 6.02 */
/*   on Wed Mar 15 14:30:09 2017 */

import functions::*;
import types::*;
import parameters::*;

/* FPGA module FM-XC7V2000T-R2 */
module mb_1_TA1 (
    clk0_p,
    clk0_n,

    sync0_p,
    sync0_n,

    dmbi_h2f,
    dmbi_f2h,

    clk1_p,
    clk1_n,

    sync1_p,
    sync1_n,

    led_red,
    led_green,
    led_blue,
    led_yellow,

    `ifdef EN_DDR
        clk2_p,
        clk2_n,
    `endif

    // SSRAM interface
    sram0_k_p,
    sram0_k_n,
    sram0_a,
    sram0_dq,
    sram0_bws_n,
    sram0_rnw,
    sram0_ld_n,
    sram0_doff_n,

    sram1_k_p,
    sram1_k_n,
    sram1_a,
    sram1_dq,
    sram1_bws_n,
    sram1_rnw,
    sram1_ld_n,
    sram1_doff_n,

    sram2_k_p,
    sram2_k_n,
    sram2_a,
    sram2_dq,
    sram2_bws_n,
    sram2_rnw,
    sram2_ld_n,
    sram2_doff_n,

    sram3_k_p,
    sram3_k_n,
    sram3_a,
    sram3_dq,
    sram3_bws_n,
    sram3_rnw,
    sram3_ld_n,
    sram3_doff_n,

    `ifdef EN_DDR
        ddr3_dq,
        ddr3_dqs_p,
        ddr3_dqs_n,
        ddr3_addr,
        ddr3_ba ,
        ddr3_ras_n,
        ddr3_cas_n ,
        ddr3_we_n   ,
        ddr3_reset_n,
        ddr3_ck_p,
        ddr3_ck_n,
        ddr3_cke ,
        ddr3_cs_n ,
        ddr3_dm ,
        ddr3_odt,
    `endif

    `ifdef EN_ETH
        eth_clk_to_mac,
        eth_col_clk_mac_freq,
        eth_crs_rgmii_sel0,
        eth_gtx_clk_tck,
        eth_mdc,
        eth_mdio,
        eth_ninterrupt,
        eth_nreset,
        eth_rx_clk,
        eth_rx_dv_rck,
        eth_rx_er_rxdv_er,
        eth_rxd,
        eth_tx_clk_rgmii_sel1,
        eth_tx_en_txen_er,
        eth_tx_er,
        eth_txd,
    `endif

    mb1_BA1_CLKIO_N_0_mb1_BC1_CLKIO_N_7,  /* BA1_CLKIO_N_0 */
    mb1_BA1_CLKIO_N_1_mb1_BC1_CLKIO_N_6,  /* BA1_CLKIO_N_1 */
    mb1_BA1_CLKIO_N_2_mb1_BC1_CLKIO_N_4,  /* BA1_CLKIO_N_2 */
    mb1_BA1_CLKIO_N_3_mb1_BC1_CLKIO_N_3,  /* BA1_CLKIO_N_3 */
    mb1_BA1_CLKIO_N_4_mb1_BC1_CLKIO_N_2,  /* BA1_CLKIO_N_4 */
    mb1_BA1_CLKIO_N_5_mb1_BC1_IO_010,  /* BA1_CLKIO_N_5 */
    mb1_BA1_CLKIO_N_6_mb1_BC1_CLKIO_N_1,  /* BA1_CLKIO_N_6 */
    mb1_BA1_CLKIO_N_7_mb1_BC1_CLKIO_N_0,  /* BA1_CLKIO_N_7 */
    mb1_BA1_CLKIO_P_0_mb1_BC1_CLKIO_P_7,  /* BA1_CLKIO_P_0 */
    mb1_BA1_CLKIO_P_1_mb1_BC1_CLKIO_P_6,  /* BA1_CLKIO_P_1 */
    mb1_BA1_CLKIO_P_2_mb1_BC1_CLKIO_P_4,  /* BA1_CLKIO_P_2 */
    mb1_BA1_CLKIO_P_3_mb1_BC1_CLKIO_P_3,  /* BA1_CLKIO_P_3 */
    mb1_BA1_CLKIO_P_4_mb1_BC1_CLKIO_P_2,  /* BA1_CLKIO_P_4 */
    mb1_BA1_CLKIO_P_5_mb1_BC1_IO_011,  /* BA1_CLKIO_P_5 */
    mb1_BA1_CLKIO_P_6_mb1_BC1_CLKIO_P_1,  /* BA1_CLKIO_P_6 */
    mb1_BA1_CLKIO_P_7_mb1_BC1_CLKIO_P_0,  /* BA1_CLKIO_P_7 */
    mb1_BA1_IO_004_mb1_BC1_IO_006,  /* BA1_IO_004 */
    mb1_BA1_IO_005_mb1_BC1_IO_007,  /* BA1_IO_005 */
    mb1_BA1_IO_006_mb1_BC1_IO_004,  /* BA1_IO_006 */
    mb1_BA1_IO_007_mb1_BC1_IO_005,  /* BA1_IO_007 */
    mb1_BA1_IO_008_mb1_BC1_IO_022,  /* BA1_IO_008 */
    mb1_BA1_IO_009_mb1_BC1_IO_023,  /* BA1_IO_009 */
    mb1_BA1_IO_010_mb1_BC1_CLKIO_N_5,  /* BA1_IO_010 */
    mb1_BA1_IO_011_mb1_BC1_CLKIO_P_5,  /* BA1_IO_011 */
    mb1_BA1_IO_012_mb1_BC1_IO_012,  /* BA1_IO_012 */
    mb1_BA1_IO_013_mb1_BC1_IO_013,  /* BA1_IO_013 */
    mb1_BA1_IO_014_mb1_BC1_IO_016,  /* BA1_IO_014 */
    mb1_BA1_IO_015_mb1_BC1_IO_017,  /* BA1_IO_015 */
    mb1_BA1_IO_016_mb1_BC1_IO_014,  /* BA1_IO_016 */
    mb1_BA1_IO_017_mb1_BC1_IO_015,  /* BA1_IO_017 */
    mb1_BA1_IO_018_mb1_BC1_IO_032,  /* BA1_IO_018 */
    mb1_BA1_IO_019_mb1_BC1_IO_033,  /* BA1_IO_019 */
    mb1_BA1_IO_020_mb1_BC1_IO_030,  /* BA1_IO_020 */
    mb1_BA1_IO_021_mb1_BC1_IO_031,  /* BA1_IO_021 */
    mb1_BA1_IO_022_mb1_BC1_IO_008,  /* BA1_IO_022 */
    mb1_BA1_IO_023_mb1_BC1_IO_009,  /* BA1_IO_023 */
    mb1_BA1_IO_024_mb1_BC1_IO_026,  /* BA1_IO_024 */
    mb1_BA1_IO_025_mb1_BC1_IO_027,  /* BA1_IO_025 */
    mb1_BA1_IO_026_mb1_BC1_IO_024,  /* BA1_IO_026 */
    mb1_BA1_IO_027_mb1_BC1_IO_025,  /* BA1_IO_027 */
    mb1_BA1_IO_028_mb1_BC1_IO_042,  /* BA1_IO_028 */
    mb1_BA1_IO_029_mb1_BC1_IO_043,  /* BA1_IO_029 */
    mb1_BA1_IO_030_mb1_BC1_IO_020,  /* BA1_IO_030 */
    mb1_BA1_IO_031_mb1_BC1_IO_021,  /* BA1_IO_031 */
    mb1_BA1_IO_032_mb1_BC1_IO_018,  /* BA1_IO_032 */
    mb1_BA1_IO_033_mb1_BC1_IO_019,  /* BA1_IO_033 */
    mb1_BA1_IO_034_mb1_BC1_IO_036,  /* BA1_IO_034 */
    mb1_BA1_IO_035_mb1_BC1_IO_037,  /* BA1_IO_035 */
    mb1_BA1_IO_036_mb1_BC1_IO_034,  /* BA1_IO_036 */
    mb1_BA1_IO_037_mb1_BC1_IO_035,  /* BA1_IO_037 */
    mb1_BA1_IO_038_mb1_BC1_IO_052,  /* BA1_IO_038 */
    mb1_BA1_IO_039_mb1_BC1_IO_053,  /* BA1_IO_039 */
    mb1_BA1_IO_040_mb1_BC1_IO_050,  /* BA1_IO_040 */
    mb1_BA1_IO_041_mb1_BC1_IO_051,  /* BA1_IO_041 */
    mb1_BA1_IO_042_mb1_BC1_IO_028,  /* BA1_IO_042 */
    mb1_BA1_IO_043_mb1_BC1_IO_029,  /* BA1_IO_043 */
    mb1_BA1_IO_044_mb1_BC1_IO_046,  /* BA1_IO_044 */
    mb1_BA1_IO_045_mb1_BC1_IO_047,  /* BA1_IO_045 */
    mb1_BA1_IO_046_mb1_BC1_IO_044,  /* BA1_IO_046 */
    mb1_BA1_IO_047_mb1_BC1_IO_045,  /* BA1_IO_047 */
    mb1_BA1_IO_048_mb1_BC1_IO_062,  /* BA1_IO_048 */
    mb1_BA1_IO_049_mb1_BC1_IO_063,  /* BA1_IO_049 */
    mb1_BA1_IO_050_mb1_BC1_IO_040,  /* BA1_IO_050 */
    mb1_BA1_IO_051_mb1_BC1_IO_041,  /* BA1_IO_051 */
    mb1_BA1_IO_052_mb1_BC1_IO_038,  /* BA1_IO_052 */
    mb1_BA1_IO_053_mb1_BC1_IO_039,  /* BA1_IO_053 */
    mb1_BA1_IO_054_mb1_BC1_IO_056,  /* BA1_IO_054 */
    mb1_BA1_IO_055_mb1_BC1_IO_057,  /* BA1_IO_055 */
    mb1_BA1_IO_056_mb1_BC1_IO_054,  /* BA1_IO_056 */
    mb1_BA1_IO_057_mb1_BC1_IO_055,  /* BA1_IO_057 */
    mb1_BA1_IO_058_mb1_BC1_IO_072,  /* BA1_IO_058 */
    mb1_BA1_IO_059_mb1_BC1_IO_073,  /* BA1_IO_059 */
    mb1_BA1_IO_060_mb1_BC1_IO_070,  /* BA1_IO_060 */
    mb1_BA1_IO_061_mb1_BC1_IO_071,  /* BA1_IO_061 */
    mb1_BA1_IO_062_mb1_BC1_IO_048,  /* BA1_IO_062 */
    mb1_BA1_IO_063_mb1_BC1_IO_049,  /* BA1_IO_063 */
    mb1_BA1_IO_064_mb1_BC1_IO_066,  /* BA1_IO_064 */
    mb1_BA1_IO_065_mb1_BC1_IO_067,  /* BA1_IO_065 */
    mb1_BA1_IO_066_mb1_BC1_IO_064,  /* BA1_IO_066 */
    mb1_BA1_IO_067_mb1_BC1_IO_065,  /* BA1_IO_067 */
    mb1_BA1_IO_068_mb1_BC1_IO_082,  /* BA1_IO_068 */
    mb1_BA1_IO_069_mb1_BC1_IO_083,  /* BA1_IO_069 */
    mb1_BA1_IO_070_mb1_BC1_IO_060,  /* BA1_IO_070 */
    mb1_BA1_IO_071_mb1_BC1_IO_061,  /* BA1_IO_071 */
    mb1_BA1_IO_072_mb1_BC1_IO_058,  /* BA1_IO_072 */
    mb1_BA1_IO_073_mb1_BC1_IO_059,  /* BA1_IO_073 */
    mb1_BA1_IO_074_mb1_BC1_IO_076,  /* BA1_IO_074 */
    mb1_BA1_IO_075_mb1_BC1_IO_077,  /* BA1_IO_075 */
    mb1_BA1_IO_076_mb1_BC1_IO_074,  /* BA1_IO_076 */
    mb1_BA1_IO_077_mb1_BC1_IO_075,  /* BA1_IO_077 */
    mb1_BA1_IO_078_mb1_BC1_IO_092,  /* BA1_IO_078 */
    mb1_BA1_IO_079_mb1_BC1_IO_093,  /* BA1_IO_079 */
    mb1_BA1_IO_080_mb1_BC1_IO_090,  /* BA1_IO_080 */
    mb1_BA1_IO_081_mb1_BC1_IO_091,  /* BA1_IO_081 */
    mb1_BA1_IO_082_mb1_BC1_IO_068,  /* BA1_IO_082 */
    mb1_BA1_IO_083_mb1_BC1_IO_069,  /* BA1_IO_083 */
    mb1_BA1_IO_084_mb1_BC1_IO_086,  /* BA1_IO_084 */
    mb1_BA1_IO_085_mb1_BC1_IO_087,  /* BA1_IO_085 */
    mb1_BA1_IO_086_mb1_BC1_IO_084,  /* BA1_IO_086 */
    mb1_BA1_IO_087_mb1_BC1_IO_085,  /* BA1_IO_087 */
    mb1_BA1_IO_088_mb1_BC1_IO_102,  /* BA1_IO_088 */
    mb1_BA1_IO_089_mb1_BC1_IO_103,  /* BA1_IO_089 */
    mb1_BA1_IO_090_mb1_BC1_IO_080,  /* BA1_IO_090 */
    mb1_BA1_IO_091_mb1_BC1_IO_081,  /* BA1_IO_091 */
    mb1_BA1_IO_092_mb1_BC1_IO_078,  /* BA1_IO_092 */
    mb1_BA1_IO_093_mb1_BC1_IO_079,  /* BA1_IO_093 */
    mb1_BA1_IO_094_mb1_BC1_IO_096,  /* BA1_IO_094 */
    mb1_BA1_IO_095_mb1_BC1_IO_097,  /* BA1_IO_095 */
    mb1_BA1_IO_096_mb1_BC1_IO_094,  /* BA1_IO_096 */
    mb1_BA1_IO_097_mb1_BC1_IO_095,  /* BA1_IO_097 */
    mb1_BA1_IO_098_mb1_BC1_IO_112,  /* BA1_IO_098 */
    mb1_BA1_IO_099_mb1_BC1_IO_113,  /* BA1_IO_099 */
    mb1_BA1_IO_100_mb1_BC1_IO_110,  /* BA1_IO_100 */
    mb1_BA1_IO_101_mb1_BC1_IO_111,  /* BA1_IO_101 */
    mb1_BA1_IO_102_mb1_BC1_IO_088,  /* BA1_IO_102 */
    mb1_BA1_IO_103_mb1_BC1_IO_089,  /* BA1_IO_103 */
    mb1_BA1_IO_104_mb1_BC1_IO_106,  /* BA1_IO_104 */
    mb1_BA1_IO_105_mb1_BC1_IO_107,  /* BA1_IO_105 */

    mb1_BB1_CLKIO_N_0_mb1_BB3_CLKIO_N_7,  /* BB1_CLKIO_N_0 */
    mb1_BB1_CLKIO_N_1_mb1_BB3_CLKIO_N_6,  /* BB1_CLKIO_N_1 */
    mb1_BB1_CLKIO_N_2_mb1_BB3_CLKIO_N_4,  /* BB1_CLKIO_N_2 */
    mb1_BB1_CLKIO_N_3_mb1_BB3_CLKIO_N_3,  /* BB1_CLKIO_N_3 */
    mb1_BB1_CLKIO_N_4_mb1_BB3_CLKIO_N_2,  /* BB1_CLKIO_N_4 */
    mb1_BB1_CLKIO_N_5_mb1_BB3_IO_010,  /* BB1_CLKIO_N_5 */
    mb1_BB1_CLKIO_N_6_mb1_BB3_CLKIO_N_1,  /* BB1_CLKIO_N_6 */
    mb1_BB1_CLKIO_N_7_mb1_BB3_CLKIO_N_0,  /* BB1_CLKIO_N_7 */
    mb1_BB1_CLKIO_P_0_mb1_BB3_CLKIO_P_7,  /* BB1_CLKIO_P_0 */
    mb1_BB1_CLKIO_P_1_mb1_BB3_CLKIO_P_6,  /* BB1_CLKIO_P_1 */
    mb1_BB1_CLKIO_P_2_mb1_BB3_CLKIO_P_4,  /* BB1_CLKIO_P_2 */
    mb1_BB1_CLKIO_P_3_mb1_BB3_CLKIO_P_3,  /* BB1_CLKIO_P_3 */
    mb1_BB1_CLKIO_P_4_mb1_BB3_CLKIO_P_2,  /* BB1_CLKIO_P_4 */
    mb1_BB1_CLKIO_P_5_mb1_BB3_IO_011,  /* BB1_CLKIO_P_5 */
    mb1_BB1_CLKIO_P_6_mb1_BB3_CLKIO_P_1,  /* BB1_CLKIO_P_6 */
    mb1_BB1_CLKIO_P_7_mb1_BB3_CLKIO_P_0,  /* BB1_CLKIO_P_7 */
    mb1_BB1_IO_004_mb1_BB3_IO_006,  /* BB1_IO_004 */
    mb1_BB1_IO_005_mb1_BB3_IO_007,  /* BB1_IO_005 */
    mb1_BB1_IO_006_mb1_BB3_IO_004,  /* BB1_IO_006 */
    mb1_BB1_IO_007_mb1_BB3_IO_005,  /* BB1_IO_007 */
    mb1_BB1_IO_008_mb1_BB3_IO_022,  /* BB1_IO_008 */
    mb1_BB1_IO_009_mb1_BB3_IO_023,  /* BB1_IO_009 */
    mb1_BB1_IO_010_mb1_BB3_CLKIO_N_5,  /* BB1_IO_010 */
    mb1_BB1_IO_011_mb1_BB3_CLKIO_P_5,  /* BB1_IO_011 */
    mb1_BB1_IO_012_mb1_BB3_IO_012,  /* BB1_IO_012 */
    mb1_BB1_IO_013_mb1_BB3_IO_013,  /* BB1_IO_013 */
    mb1_BB1_IO_014_mb1_BB3_IO_016,  /* BB1_IO_014 */
    mb1_BB1_IO_015_mb1_BB3_IO_017,  /* BB1_IO_015 */
    mb1_BB1_IO_016_mb1_BB3_IO_014,  /* BB1_IO_016 */
    mb1_BB1_IO_017_mb1_BB3_IO_015,  /* BB1_IO_017 */
    mb1_BB1_IO_018_mb1_BB3_IO_032,  /* BB1_IO_018 */
    mb1_BB1_IO_019_mb1_BB3_IO_033,  /* BB1_IO_019 */
    mb1_BB1_IO_020_mb1_BB3_IO_030,  /* BB1_IO_020 */
    mb1_BB1_IO_021_mb1_BB3_IO_031,  /* BB1_IO_021 */
    mb1_BB1_IO_022_mb1_BB3_IO_008,  /* BB1_IO_022 */
    mb1_BB1_IO_023_mb1_BB3_IO_009,  /* BB1_IO_023 */
    mb1_BB1_IO_024_mb1_BB3_IO_026,  /* BB1_IO_024 */
    mb1_BB1_IO_025_mb1_BB3_IO_027,  /* BB1_IO_025 */
    mb1_BB1_IO_026_mb1_BB3_IO_024,  /* BB1_IO_026 */
    mb1_BB1_IO_027_mb1_BB3_IO_025,  /* BB1_IO_027 */
    mb1_BB1_IO_028_mb1_BB3_IO_042,  /* BB1_IO_028 */
    mb1_BB1_IO_029_mb1_BB3_IO_043,  /* BB1_IO_029 */
    mb1_BB1_IO_030_mb1_BB3_IO_020,  /* BB1_IO_030 */
    mb1_BB1_IO_031_mb1_BB3_IO_021,  /* BB1_IO_031 */
    mb1_BB1_IO_032_mb1_BB3_IO_018,  /* BB1_IO_032 */
    mb1_BB1_IO_033_mb1_BB3_IO_019,  /* BB1_IO_033 */
    mb1_BB1_IO_034_mb1_BB3_IO_036,  /* BB1_IO_034 */
    mb1_BB1_IO_035_mb1_BB3_IO_037,  /* BB1_IO_035 */
    mb1_BB1_IO_036_mb1_BB3_IO_034,  /* BB1_IO_036 */
    mb1_BB1_IO_037_mb1_BB3_IO_035,  /* BB1_IO_037 */
    mb1_BB1_IO_038_mb1_BB3_IO_052,  /* BB1_IO_038 */
    mb1_BB1_IO_039_mb1_BB3_IO_053,  /* BB1_IO_039 */
    mb1_BB1_IO_040_mb1_BB3_IO_050,  /* BB1_IO_040 */
    mb1_BB1_IO_041_mb1_BB3_IO_051,  /* BB1_IO_041 */
    mb1_BB1_IO_042_mb1_BB3_IO_028,  /* BB1_IO_042 */
    mb1_BB1_IO_043_mb1_BB3_IO_029,  /* BB1_IO_043 */
    mb1_BB1_IO_044_mb1_BB3_IO_046,  /* BB1_IO_044 */
    mb1_BB1_IO_045_mb1_BB3_IO_047,  /* BB1_IO_045 */
    mb1_BB1_IO_046_mb1_BB3_IO_044,  /* BB1_IO_046 */
    mb1_BB1_IO_047_mb1_BB3_IO_045,  /* BB1_IO_047 */
    mb1_BB1_IO_048_mb1_BB3_IO_062,  /* BB1_IO_048 */
    mb1_BB1_IO_049_mb1_BB3_IO_063,  /* BB1_IO_049 */
    mb1_BB1_IO_050_mb1_BB3_IO_040,  /* BB1_IO_050 */
    mb1_BB1_IO_051_mb1_BB3_IO_041,  /* BB1_IO_051 */
    mb1_BB1_IO_052_mb1_BB3_IO_038,  /* BB1_IO_052 */
    mb1_BB1_IO_053_mb1_BB3_IO_039,  /* BB1_IO_053 */
    mb1_BB1_IO_054_mb1_BB3_IO_056,  /* BB1_IO_054 */
    mb1_BB1_IO_055_mb1_BB3_IO_057,  /* BB1_IO_055 */
    mb1_BB1_IO_056_mb1_BB3_IO_054,  /* BB1_IO_056 */
    mb1_BB1_IO_057_mb1_BB3_IO_055,  /* BB1_IO_057 */
    mb1_BB1_IO_058_mb1_BB3_IO_072,  /* BB1_IO_058 */
    mb1_BB1_IO_059_mb1_BB3_IO_073,  /* BB1_IO_059 */
    mb1_BB1_IO_060_mb1_BB3_IO_070,  /* BB1_IO_060 */
    mb1_BB1_IO_061_mb1_BB3_IO_071,  /* BB1_IO_061 */
    mb1_BB1_IO_062_mb1_BB3_IO_048,  /* BB1_IO_062 */
    mb1_BB1_IO_063_mb1_BB3_IO_049,  /* BB1_IO_063 */
    mb1_BB1_IO_064_mb1_BB3_IO_066,  /* BB1_IO_064 */
    mb1_BB1_IO_065_mb1_BB3_IO_067,  /* BB1_IO_065 */
    mb1_BB1_IO_066_mb1_BB3_IO_064,  /* BB1_IO_066 */
    mb1_BB1_IO_067_mb1_BB3_IO_065,  /* BB1_IO_067 */
    mb1_BB1_IO_068_mb1_BB3_IO_082,  /* BB1_IO_068 */
    mb1_BB1_IO_069_mb1_BB3_IO_083,  /* BB1_IO_069 */
    mb1_BB1_IO_070_mb1_BB3_IO_060,  /* BB1_IO_070 */
    mb1_BB1_IO_071_mb1_BB3_IO_061,  /* BB1_IO_071 */
    mb1_BB1_IO_072_mb1_BB3_IO_058,  /* BB1_IO_072 */
    mb1_BB1_IO_073_mb1_BB3_IO_059,  /* BB1_IO_073 */
    mb1_BB1_IO_074_mb1_BB3_IO_076,  /* BB1_IO_074 */
    mb1_BB1_IO_075_mb1_BB3_IO_077,  /* BB1_IO_075 */
    mb1_BB1_IO_076_mb1_BB3_IO_074,  /* BB1_IO_076 */
    mb1_BB1_IO_077_mb1_BB3_IO_075,  /* BB1_IO_077 */
    mb1_BB1_IO_078_mb1_BB3_IO_092,  /* BB1_IO_078 */
    mb1_BB1_IO_079_mb1_BB3_IO_093,  /* BB1_IO_079 */
    mb1_BB1_IO_080_mb1_BB3_IO_090,  /* BB1_IO_080 */
    mb1_BB1_IO_081_mb1_BB3_IO_091,  /* BB1_IO_081 */
    mb1_BB1_IO_082_mb1_BB3_IO_068,  /* BB1_IO_082 */
    mb1_BB1_IO_083_mb1_BB3_IO_069,  /* BB1_IO_083 */
    mb1_BB1_IO_084_mb1_BB3_IO_086,  /* BB1_IO_084 */
    mb1_BB1_IO_085_mb1_BB3_IO_087,  /* BB1_IO_085 */
    mb1_BB1_IO_086_mb1_BB3_IO_084,  /* BB1_IO_086 */
    mb1_BB1_IO_087_mb1_BB3_IO_085,  /* BB1_IO_087 */
    mb1_BB1_IO_088_mb1_BB3_IO_102,  /* BB1_IO_088 */
    mb1_BB1_IO_089_mb1_BB3_IO_103,  /* BB1_IO_089 */
    mb1_BB1_IO_090_mb1_BB3_IO_080,  /* BB1_IO_090 */
    mb1_BB1_IO_091_mb1_BB3_IO_081,  /* BB1_IO_091 */
    mb1_BB1_IO_092_mb1_BB3_IO_078,  /* BB1_IO_092 */
    mb1_BB1_IO_093_mb1_BB3_IO_079,  /* BB1_IO_093 */
    mb1_BB1_IO_094_mb1_BB3_IO_096,  /* BB1_IO_094 */
    mb1_BB1_IO_095_mb1_BB3_IO_097,  /* BB1_IO_095 */
    mb1_BB1_IO_096_mb1_BB3_IO_094,  /* BB1_IO_096 */
    mb1_BB1_IO_097_mb1_BB3_IO_095,  /* BB1_IO_097 */
    mb1_BB1_IO_098_mb1_BB3_IO_112,  /* BB1_IO_098 */
    mb1_BB1_IO_099_mb1_BB3_IO_113,  /* BB1_IO_099 */
    mb1_BB1_IO_100_mb1_BB3_IO_110,  /* BB1_IO_100 */
    mb1_BB1_IO_101_mb1_BB3_IO_111,  /* BB1_IO_101 */
    mb1_BB1_IO_102_mb1_BB3_IO_088,  /* BB1_IO_102 */
    mb1_BB1_IO_103_mb1_BB3_IO_089,  /* BB1_IO_103 */
    mb1_BB1_IO_104_mb1_BB3_IO_106,  /* BB1_IO_104 */
    mb1_BB1_IO_105_mb1_BB3_IO_107   /* BB1_IO_105 */
    );

    /* pins which are not connected to an x-board */
    parameter ADDR_W  = 22;
    parameter DQ_PINS = 18;
    parameter GROUPS  = 2;

    output logic               sram0_k_p;
    output logic               sram0_k_n;
    output logic [ADDR_W-1:0]  sram0_a;
    inout  tri   [DQ_PINS-1:0] sram0_dq;
    output logic [GROUPS-1:0]  sram0_bws_n;
    output logic               sram0_rnw;
    output logic               sram0_ld_n;
    output logic               sram0_doff_n;

    output logic               sram1_k_p;
    output logic               sram1_k_n;
    output logic [ADDR_W-1:0]  sram1_a;
    inout  tri   [DQ_PINS-1:0] sram1_dq;
    output logic [GROUPS-1:0]  sram1_bws_n;
    output logic               sram1_rnw;
    output logic               sram1_ld_n;
    output logic               sram1_doff_n;

    output logic               sram2_k_p;
    output logic               sram2_k_n;
    output logic [ADDR_W-1:0]  sram2_a;
    inout  tri   [DQ_PINS-1:0] sram2_dq;
    output logic [GROUPS-1:0]  sram2_bws_n;
    output logic               sram2_rnw;
    output logic               sram2_ld_n;
    output logic               sram2_doff_n;

    output logic               sram3_k_p;
    output logic               sram3_k_n;
    output logic [ADDR_W-1:0]  sram3_a;
    inout  tri   [DQ_PINS-1:0] sram3_dq;
    output logic [GROUPS-1:0]  sram3_bws_n;
    output logic               sram3_rnw;
    output logic               sram3_ld_n;
    output logic               sram3_doff_n;

    `ifdef EN_DDR
        inout wire  [63:0] ddr3_dq;
        inout wire  [7:0]  ddr3_dqs_n;
        inout wire  [7:0]  ddr3_dqs_p;
        output wire [14:0] ddr3_addr;
        output wire [2:0]  ddr3_ba;
        output wire        ddr3_ras_n;
        output wire        ddr3_cas_n;
        output wire        ddr3_we_n;
        output wire        ddr3_reset_n;
        output wire        ddr3_ck_p;
        output wire        ddr3_ck_n;
        output wire        ddr3_cke;
        output wire        ddr3_cs_n;
        output wire [7:0]  ddr3_dm;
        output wire        ddr3_odt;
    `endif

    `ifdef EN_ETH
        input  logic       eth_clk_to_mac;
        input  logic       eth_col_clk_mac_freq;
        input  logic       eth_crs_rgmii_sel0;
        output logic       eth_gtx_clk_tck;
        output logic       eth_mdc;
        inout  tri         eth_mdio;
        input  logic       eth_ninterrupt;
        output logic       eth_nreset;
        input  logic       eth_rx_clk;
        input  logic       eth_rx_dv_rck;
        input  logic       eth_rx_er_rxdv_er;
        input  logic [7:0] eth_rxd;
        input  logic       eth_tx_clk_rgmii_sel1;
        output logic       eth_tx_en_txen_er;
        output logic       eth_tx_er;
        output logic [7:0] eth_txd;
    `endif

    output logic [19:0] dmbi_f2h;
    input  logic [19:0] dmbi_h2f;

    input logic clk0_p;
    input logic clk0_n;
    input logic sync0_p;
    input logic sync0_n;

    input logic clk1_p;
    input logic clk1_n;
    input logic sync1_p;
    input logic sync1_n;

    output logic led_red;
    output logic led_green;
    output logic led_blue;
    output logic led_yellow;

    `ifdef EN_DDR
        input logic clk2_n;
        input logic clk2_p;
    `endif

    /* pins which are connected to motherboard connector BA1 */
    /* and connector BA2 on x-board IC-PDS-CABLE-R1 */
    input wire mb1_BA1_CLKIO_N_0_mb1_BC1_CLKIO_N_7;
    input wire mb1_BA1_CLKIO_N_1_mb1_BC1_CLKIO_N_6;
    input wire mb1_BA1_CLKIO_N_2_mb1_BC1_CLKIO_N_4;
    input wire mb1_BA1_CLKIO_N_3_mb1_BC1_CLKIO_N_3;
    input wire mb1_BA1_CLKIO_N_4_mb1_BC1_CLKIO_N_2;
    input wire mb1_BA1_CLKIO_N_5_mb1_BC1_IO_010;
    input wire mb1_BA1_CLKIO_N_6_mb1_BC1_CLKIO_N_1;
    input wire mb1_BA1_CLKIO_N_7_mb1_BC1_CLKIO_N_0;
    input wire mb1_BA1_CLKIO_P_0_mb1_BC1_CLKIO_P_7;
    input wire mb1_BA1_CLKIO_P_1_mb1_BC1_CLKIO_P_6;
    input wire mb1_BA1_CLKIO_P_2_mb1_BC1_CLKIO_P_4;
    input wire mb1_BA1_CLKIO_P_3_mb1_BC1_CLKIO_P_3;
    input wire mb1_BA1_CLKIO_P_4_mb1_BC1_CLKIO_P_2;
    input wire mb1_BA1_CLKIO_P_5_mb1_BC1_IO_011;
    input wire mb1_BA1_CLKIO_P_6_mb1_BC1_CLKIO_P_1;
    input wire mb1_BA1_CLKIO_P_7_mb1_BC1_CLKIO_P_0;
    input wire mb1_BA1_IO_004_mb1_BC1_IO_006;
    input wire mb1_BA1_IO_005_mb1_BC1_IO_007;
    input wire mb1_BA1_IO_006_mb1_BC1_IO_004;
    input wire mb1_BA1_IO_007_mb1_BC1_IO_005;
    input wire mb1_BA1_IO_008_mb1_BC1_IO_022;
    input wire mb1_BA1_IO_009_mb1_BC1_IO_023;
    input wire mb1_BA1_IO_010_mb1_BC1_CLKIO_N_5;
    input wire mb1_BA1_IO_011_mb1_BC1_CLKIO_P_5;
    input wire mb1_BA1_IO_012_mb1_BC1_IO_012;
    input wire mb1_BA1_IO_013_mb1_BC1_IO_013;
    input wire mb1_BA1_IO_014_mb1_BC1_IO_016;
    input wire mb1_BA1_IO_015_mb1_BC1_IO_017;
    input wire mb1_BA1_IO_016_mb1_BC1_IO_014;
    input wire mb1_BA1_IO_017_mb1_BC1_IO_015;
    input wire mb1_BA1_IO_018_mb1_BC1_IO_032;
    input wire mb1_BA1_IO_019_mb1_BC1_IO_033;
    input wire mb1_BA1_IO_020_mb1_BC1_IO_030;
    input wire mb1_BA1_IO_021_mb1_BC1_IO_031;
    input wire mb1_BA1_IO_022_mb1_BC1_IO_008;
    input wire mb1_BA1_IO_023_mb1_BC1_IO_009;
    input wire mb1_BA1_IO_024_mb1_BC1_IO_026;
    input wire mb1_BA1_IO_025_mb1_BC1_IO_027;
    input wire mb1_BA1_IO_026_mb1_BC1_IO_024;
    input wire mb1_BA1_IO_027_mb1_BC1_IO_025;
    input wire mb1_BA1_IO_028_mb1_BC1_IO_042;
    input wire mb1_BA1_IO_029_mb1_BC1_IO_043;
    input wire mb1_BA1_IO_030_mb1_BC1_IO_020;
    input wire mb1_BA1_IO_031_mb1_BC1_IO_021;
    input wire mb1_BA1_IO_032_mb1_BC1_IO_018;
    input wire mb1_BA1_IO_033_mb1_BC1_IO_019;
    input wire mb1_BA1_IO_034_mb1_BC1_IO_036;
    input wire mb1_BA1_IO_035_mb1_BC1_IO_037;
    input wire mb1_BA1_IO_036_mb1_BC1_IO_034;
    input wire mb1_BA1_IO_037_mb1_BC1_IO_035;
    input wire mb1_BA1_IO_038_mb1_BC1_IO_052;
    input wire mb1_BA1_IO_039_mb1_BC1_IO_053;
    input wire mb1_BA1_IO_040_mb1_BC1_IO_050;
    input wire mb1_BA1_IO_041_mb1_BC1_IO_051;
    input wire mb1_BA1_IO_042_mb1_BC1_IO_028;
    input wire mb1_BA1_IO_043_mb1_BC1_IO_029;
    input wire mb1_BA1_IO_044_mb1_BC1_IO_046;
    input wire mb1_BA1_IO_045_mb1_BC1_IO_047;
    input wire mb1_BA1_IO_046_mb1_BC1_IO_044;
    output wire mb1_BA1_IO_047_mb1_BC1_IO_045;
    output wire mb1_BA1_IO_048_mb1_BC1_IO_062;
    output wire mb1_BA1_IO_049_mb1_BC1_IO_063;
    output wire mb1_BA1_IO_050_mb1_BC1_IO_040;
    output wire mb1_BA1_IO_051_mb1_BC1_IO_041;
    output wire mb1_BA1_IO_052_mb1_BC1_IO_038;
    output wire mb1_BA1_IO_053_mb1_BC1_IO_039;
    output wire mb1_BA1_IO_054_mb1_BC1_IO_056;
    output wire mb1_BA1_IO_055_mb1_BC1_IO_057;
    output wire mb1_BA1_IO_056_mb1_BC1_IO_054;
    output wire mb1_BA1_IO_057_mb1_BC1_IO_055;
    output wire mb1_BA1_IO_058_mb1_BC1_IO_072;
    output wire mb1_BA1_IO_059_mb1_BC1_IO_073;
    output wire mb1_BA1_IO_060_mb1_BC1_IO_070;
    output wire mb1_BA1_IO_061_mb1_BC1_IO_071;
    output wire mb1_BA1_IO_062_mb1_BC1_IO_048;
    output wire mb1_BA1_IO_063_mb1_BC1_IO_049;
    output wire mb1_BA1_IO_064_mb1_BC1_IO_066;
    output wire mb1_BA1_IO_065_mb1_BC1_IO_067;
    output wire mb1_BA1_IO_066_mb1_BC1_IO_064;
    output wire mb1_BA1_IO_067_mb1_BC1_IO_065;
    output wire mb1_BA1_IO_068_mb1_BC1_IO_082;
    output wire mb1_BA1_IO_069_mb1_BC1_IO_083;
    output wire mb1_BA1_IO_070_mb1_BC1_IO_060;
    output wire mb1_BA1_IO_071_mb1_BC1_IO_061;
    output wire mb1_BA1_IO_072_mb1_BC1_IO_058;
    output wire mb1_BA1_IO_073_mb1_BC1_IO_059;
    output wire mb1_BA1_IO_074_mb1_BC1_IO_076;
    output wire mb1_BA1_IO_075_mb1_BC1_IO_077;
    output wire mb1_BA1_IO_076_mb1_BC1_IO_074;
    output wire mb1_BA1_IO_077_mb1_BC1_IO_075;
    output wire mb1_BA1_IO_078_mb1_BC1_IO_092;
    output wire mb1_BA1_IO_079_mb1_BC1_IO_093;
    output wire mb1_BA1_IO_080_mb1_BC1_IO_090;
    output wire mb1_BA1_IO_081_mb1_BC1_IO_091;
    output wire mb1_BA1_IO_082_mb1_BC1_IO_068;
    output wire mb1_BA1_IO_083_mb1_BC1_IO_069;
    output wire mb1_BA1_IO_084_mb1_BC1_IO_086;
    output wire mb1_BA1_IO_085_mb1_BC1_IO_087;
    output wire mb1_BA1_IO_086_mb1_BC1_IO_084;
    output wire mb1_BA1_IO_087_mb1_BC1_IO_085;
    output wire mb1_BA1_IO_088_mb1_BC1_IO_102;
    output wire mb1_BA1_IO_089_mb1_BC1_IO_103;
    output wire mb1_BA1_IO_090_mb1_BC1_IO_080;
    output wire mb1_BA1_IO_091_mb1_BC1_IO_081;
    output wire mb1_BA1_IO_092_mb1_BC1_IO_078;
    output wire mb1_BA1_IO_093_mb1_BC1_IO_079;
    output wire mb1_BA1_IO_094_mb1_BC1_IO_096;
    output wire mb1_BA1_IO_095_mb1_BC1_IO_097;
    output wire mb1_BA1_IO_096_mb1_BC1_IO_094;
    output wire mb1_BA1_IO_097_mb1_BC1_IO_095;
    output wire mb1_BA1_IO_098_mb1_BC1_IO_112;
    output wire mb1_BA1_IO_099_mb1_BC1_IO_113;
    output wire mb1_BA1_IO_100_mb1_BC1_IO_110;
    output wire mb1_BA1_IO_101_mb1_BC1_IO_111;
    output wire mb1_BA1_IO_102_mb1_BC1_IO_088;
    output wire mb1_BA1_IO_103_mb1_BC1_IO_089;
    output wire mb1_BA1_IO_104_mb1_BC1_IO_106;
    output wire mb1_BA1_IO_105_mb1_BC1_IO_107;

    /* pins which are connected to motherboard connector BB1 */
    /* and connector BA1 on x-board IC-PDS-CABLE-R1 */
    input wire mb1_BB1_CLKIO_N_0_mb1_BB3_CLKIO_N_7;
    input wire mb1_BB1_CLKIO_N_1_mb1_BB3_CLKIO_N_6;
    input wire mb1_BB1_CLKIO_N_2_mb1_BB3_CLKIO_N_4;
    input wire mb1_BB1_CLKIO_N_3_mb1_BB3_CLKIO_N_3;
    input wire mb1_BB1_CLKIO_N_4_mb1_BB3_CLKIO_N_2;
    input wire mb1_BB1_CLKIO_N_5_mb1_BB3_IO_010;
    input wire mb1_BB1_CLKIO_N_6_mb1_BB3_CLKIO_N_1;
    input wire mb1_BB1_CLKIO_N_7_mb1_BB3_CLKIO_N_0;
    input wire mb1_BB1_CLKIO_P_0_mb1_BB3_CLKIO_P_7;
    input wire mb1_BB1_CLKIO_P_1_mb1_BB3_CLKIO_P_6;
    input wire mb1_BB1_CLKIO_P_2_mb1_BB3_CLKIO_P_4;
    input wire mb1_BB1_CLKIO_P_3_mb1_BB3_CLKIO_P_3;
    input wire mb1_BB1_CLKIO_P_4_mb1_BB3_CLKIO_P_2;
    input wire mb1_BB1_CLKIO_P_5_mb1_BB3_IO_011;
    input wire mb1_BB1_CLKIO_P_6_mb1_BB3_CLKIO_P_1;
    input wire mb1_BB1_CLKIO_P_7_mb1_BB3_CLKIO_P_0;
    input wire mb1_BB1_IO_004_mb1_BB3_IO_006;
    input wire mb1_BB1_IO_005_mb1_BB3_IO_007;
    input wire mb1_BB1_IO_006_mb1_BB3_IO_004;
    input wire mb1_BB1_IO_007_mb1_BB3_IO_005;
    input wire mb1_BB1_IO_008_mb1_BB3_IO_022;
    input wire mb1_BB1_IO_009_mb1_BB3_IO_023;
    input wire mb1_BB1_IO_010_mb1_BB3_CLKIO_N_5;
    input wire mb1_BB1_IO_011_mb1_BB3_CLKIO_P_5;
    input wire mb1_BB1_IO_012_mb1_BB3_IO_012;
    input wire mb1_BB1_IO_013_mb1_BB3_IO_013;
    input wire mb1_BB1_IO_014_mb1_BB3_IO_016;
    input wire mb1_BB1_IO_015_mb1_BB3_IO_017;
    input wire mb1_BB1_IO_016_mb1_BB3_IO_014;
    input wire mb1_BB1_IO_017_mb1_BB3_IO_015;
    input wire mb1_BB1_IO_018_mb1_BB3_IO_032;
    input wire mb1_BB1_IO_019_mb1_BB3_IO_033;
    input wire mb1_BB1_IO_020_mb1_BB3_IO_030;
    input wire mb1_BB1_IO_021_mb1_BB3_IO_031;
    input wire mb1_BB1_IO_022_mb1_BB3_IO_008;
    input wire mb1_BB1_IO_023_mb1_BB3_IO_009;
    input wire mb1_BB1_IO_024_mb1_BB3_IO_026;
    input wire mb1_BB1_IO_025_mb1_BB3_IO_027;
    input wire mb1_BB1_IO_026_mb1_BB3_IO_024;
    input wire mb1_BB1_IO_027_mb1_BB3_IO_025;
    input wire mb1_BB1_IO_028_mb1_BB3_IO_042;
    input wire mb1_BB1_IO_029_mb1_BB3_IO_043;
    input wire mb1_BB1_IO_030_mb1_BB3_IO_020;
    input wire mb1_BB1_IO_031_mb1_BB3_IO_021;
    input wire mb1_BB1_IO_032_mb1_BB3_IO_018;
    input wire mb1_BB1_IO_033_mb1_BB3_IO_019;
    input wire mb1_BB1_IO_034_mb1_BB3_IO_036;
    input wire mb1_BB1_IO_035_mb1_BB3_IO_037;
    input wire mb1_BB1_IO_036_mb1_BB3_IO_034;
    input wire mb1_BB1_IO_037_mb1_BB3_IO_035;
    input wire mb1_BB1_IO_038_mb1_BB3_IO_052;
    input wire mb1_BB1_IO_039_mb1_BB3_IO_053;
    input wire mb1_BB1_IO_040_mb1_BB3_IO_050;
    input wire mb1_BB1_IO_041_mb1_BB3_IO_051;
    input wire mb1_BB1_IO_042_mb1_BB3_IO_028;
    input wire mb1_BB1_IO_043_mb1_BB3_IO_029;
    input wire mb1_BB1_IO_044_mb1_BB3_IO_046;
    input wire mb1_BB1_IO_045_mb1_BB3_IO_047;
    input wire mb1_BB1_IO_046_mb1_BB3_IO_044;
    output wire mb1_BB1_IO_047_mb1_BB3_IO_045;
    output wire mb1_BB1_IO_048_mb1_BB3_IO_062;
    output wire mb1_BB1_IO_049_mb1_BB3_IO_063;
    output wire mb1_BB1_IO_050_mb1_BB3_IO_040;
    output wire mb1_BB1_IO_051_mb1_BB3_IO_041;
    output wire mb1_BB1_IO_052_mb1_BB3_IO_038;
    output wire mb1_BB1_IO_053_mb1_BB3_IO_039;
    output wire mb1_BB1_IO_054_mb1_BB3_IO_056;
    output wire mb1_BB1_IO_055_mb1_BB3_IO_057;
    output wire mb1_BB1_IO_056_mb1_BB3_IO_054;
    output wire mb1_BB1_IO_057_mb1_BB3_IO_055;
    output wire mb1_BB1_IO_058_mb1_BB3_IO_072;
    output wire mb1_BB1_IO_059_mb1_BB3_IO_073;
    output wire mb1_BB1_IO_060_mb1_BB3_IO_070;
    output wire mb1_BB1_IO_061_mb1_BB3_IO_071;
    output wire mb1_BB1_IO_062_mb1_BB3_IO_048;
    output wire mb1_BB1_IO_063_mb1_BB3_IO_049;
    output wire mb1_BB1_IO_064_mb1_BB3_IO_066;
    output wire mb1_BB1_IO_065_mb1_BB3_IO_067;
    output wire mb1_BB1_IO_066_mb1_BB3_IO_064;
    output wire mb1_BB1_IO_067_mb1_BB3_IO_065;
    output wire mb1_BB1_IO_068_mb1_BB3_IO_082;
    output wire mb1_BB1_IO_069_mb1_BB3_IO_083;
    output wire mb1_BB1_IO_070_mb1_BB3_IO_060;
    output wire mb1_BB1_IO_071_mb1_BB3_IO_061;
    output wire mb1_BB1_IO_072_mb1_BB3_IO_058;
    output wire mb1_BB1_IO_073_mb1_BB3_IO_059;
    output wire mb1_BB1_IO_074_mb1_BB3_IO_076;
    output wire mb1_BB1_IO_075_mb1_BB3_IO_077;
    output wire mb1_BB1_IO_076_mb1_BB3_IO_074;
    output wire mb1_BB1_IO_077_mb1_BB3_IO_075;
    output wire mb1_BB1_IO_078_mb1_BB3_IO_092;
    output wire mb1_BB1_IO_079_mb1_BB3_IO_093;
    output wire mb1_BB1_IO_080_mb1_BB3_IO_090;
    output wire mb1_BB1_IO_081_mb1_BB3_IO_091;
    output wire mb1_BB1_IO_082_mb1_BB3_IO_068;
    output wire mb1_BB1_IO_083_mb1_BB3_IO_069;
    output wire mb1_BB1_IO_084_mb1_BB3_IO_086;
    output wire mb1_BB1_IO_085_mb1_BB3_IO_087;
    output wire mb1_BB1_IO_086_mb1_BB3_IO_084;
    output wire mb1_BB1_IO_087_mb1_BB3_IO_085;
    output wire mb1_BB1_IO_088_mb1_BB3_IO_102;
    output wire mb1_BB1_IO_089_mb1_BB3_IO_103;
    output wire mb1_BB1_IO_090_mb1_BB3_IO_080;
    output wire mb1_BB1_IO_091_mb1_BB3_IO_081;
    output wire mb1_BB1_IO_092_mb1_BB3_IO_078;
    output wire mb1_BB1_IO_093_mb1_BB3_IO_079;
    output wire mb1_BB1_IO_094_mb1_BB3_IO_096;
    output wire mb1_BB1_IO_095_mb1_BB3_IO_097;
    output wire mb1_BB1_IO_096_mb1_BB3_IO_094;
    output wire mb1_BB1_IO_097_mb1_BB3_IO_095;
    output wire mb1_BB1_IO_098_mb1_BB3_IO_112;
    output wire mb1_BB1_IO_099_mb1_BB3_IO_113;
    output wire mb1_BB1_IO_100_mb1_BB3_IO_110;
    output wire mb1_BB1_IO_101_mb1_BB3_IO_111;
    output wire mb1_BB1_IO_102_mb1_BB3_IO_088;
    output wire mb1_BB1_IO_103_mb1_BB3_IO_089;
    output wire mb1_BB1_IO_104_mb1_BB3_IO_106;
    output wire mb1_BB1_IO_105_mb1_BB3_IO_107;

    localparam TX_PINS = 59;
    localparam RX_PINS = 59;

    wire [TX_PINS-1:0] tx_pin;
    wire [RX_PINS-1:0] rx_pin;

    assign rx_pin[0] = mb1_BA1_CLKIO_N_0_mb1_BC1_CLKIO_N_7;
    assign rx_pin[1] = mb1_BA1_CLKIO_N_1_mb1_BC1_CLKIO_N_6;
    assign rx_pin[2] = mb1_BA1_CLKIO_N_2_mb1_BC1_CLKIO_N_4;
    assign rx_pin[3] = mb1_BA1_CLKIO_N_3_mb1_BC1_CLKIO_N_3;
    assign rx_pin[4] = mb1_BA1_CLKIO_N_4_mb1_BC1_CLKIO_N_2;
    assign rx_pin[5] = mb1_BA1_CLKIO_N_5_mb1_BC1_IO_010;
    assign rx_pin[6] = mb1_BA1_CLKIO_N_6_mb1_BC1_CLKIO_N_1;
    assign rx_pin[7] = mb1_BA1_CLKIO_N_7_mb1_BC1_CLKIO_N_0;
    assign rx_pin[8] = mb1_BA1_CLKIO_P_0_mb1_BC1_CLKIO_P_7;
    assign rx_pin[9] = mb1_BA1_CLKIO_P_1_mb1_BC1_CLKIO_P_6;
    assign rx_pin[10] = mb1_BA1_CLKIO_P_2_mb1_BC1_CLKIO_P_4;
    assign rx_pin[11] = mb1_BA1_CLKIO_P_3_mb1_BC1_CLKIO_P_3;
    assign rx_pin[12] = mb1_BA1_CLKIO_P_4_mb1_BC1_CLKIO_P_2;
    assign rx_pin[13] = mb1_BA1_CLKIO_P_5_mb1_BC1_IO_011;
    assign rx_pin[14] = mb1_BA1_CLKIO_P_6_mb1_BC1_CLKIO_P_1;
    assign rx_pin[15] = mb1_BA1_CLKIO_P_7_mb1_BC1_CLKIO_P_0;
    assign rx_pin[16] = mb1_BA1_IO_004_mb1_BC1_IO_006;
    assign rx_pin[17] = mb1_BA1_IO_005_mb1_BC1_IO_007;
    assign rx_pin[18] = mb1_BA1_IO_006_mb1_BC1_IO_004;
    assign rx_pin[19] = mb1_BA1_IO_007_mb1_BC1_IO_005;
    assign rx_pin[20] = mb1_BA1_IO_008_mb1_BC1_IO_022;
    assign rx_pin[21] = mb1_BA1_IO_009_mb1_BC1_IO_023;
    assign rx_pin[22] = mb1_BA1_IO_010_mb1_BC1_CLKIO_N_5;
    assign rx_pin[23] = mb1_BA1_IO_011_mb1_BC1_CLKIO_P_5;
    assign rx_pin[24] = mb1_BA1_IO_012_mb1_BC1_IO_012;
    assign rx_pin[25] = mb1_BA1_IO_013_mb1_BC1_IO_013;
    assign rx_pin[26] = mb1_BA1_IO_014_mb1_BC1_IO_016;
    assign rx_pin[27] = mb1_BA1_IO_015_mb1_BC1_IO_017;
    assign rx_pin[28] = mb1_BA1_IO_016_mb1_BC1_IO_014;
    assign rx_pin[29] = mb1_BA1_IO_017_mb1_BC1_IO_015;
    assign rx_pin[30] = mb1_BA1_IO_018_mb1_BC1_IO_032;
    assign rx_pin[31] = mb1_BA1_IO_019_mb1_BC1_IO_033;
    assign rx_pin[32] = mb1_BA1_IO_020_mb1_BC1_IO_030;
    assign rx_pin[33] = mb1_BA1_IO_021_mb1_BC1_IO_031;
    assign rx_pin[34] = mb1_BA1_IO_022_mb1_BC1_IO_008;
    assign rx_pin[35] = mb1_BA1_IO_023_mb1_BC1_IO_009;
    assign rx_pin[36] = mb1_BA1_IO_024_mb1_BC1_IO_026;
    assign rx_pin[37] = mb1_BA1_IO_025_mb1_BC1_IO_027;
    assign rx_pin[38] = mb1_BA1_IO_026_mb1_BC1_IO_024;
    assign rx_pin[39] = mb1_BA1_IO_027_mb1_BC1_IO_025;
    assign rx_pin[40] = mb1_BA1_IO_028_mb1_BC1_IO_042;
    assign rx_pin[41] = mb1_BA1_IO_029_mb1_BC1_IO_043;
    assign rx_pin[42] = mb1_BA1_IO_030_mb1_BC1_IO_020;
    assign rx_pin[43] = mb1_BA1_IO_031_mb1_BC1_IO_021;
    assign rx_pin[44] = mb1_BA1_IO_032_mb1_BC1_IO_018;
    assign rx_pin[45] = mb1_BA1_IO_033_mb1_BC1_IO_019;
    assign rx_pin[46] = mb1_BA1_IO_034_mb1_BC1_IO_036;
    assign rx_pin[47] = mb1_BA1_IO_035_mb1_BC1_IO_037;
    assign rx_pin[48] = mb1_BA1_IO_036_mb1_BC1_IO_034;
    assign rx_pin[49] = mb1_BA1_IO_037_mb1_BC1_IO_035;
    assign rx_pin[50] = mb1_BA1_IO_038_mb1_BC1_IO_052;
    assign rx_pin[51] = mb1_BA1_IO_039_mb1_BC1_IO_053;
    assign rx_pin[52] = mb1_BA1_IO_040_mb1_BC1_IO_050;
    assign rx_pin[53] = mb1_BA1_IO_041_mb1_BC1_IO_051;
    assign rx_pin[54] = mb1_BA1_IO_042_mb1_BC1_IO_028;
    assign rx_pin[55] = mb1_BA1_IO_043_mb1_BC1_IO_029;
    assign rx_pin[56] = mb1_BA1_IO_044_mb1_BC1_IO_046;
    assign rx_pin[57] = mb1_BA1_IO_045_mb1_BC1_IO_047;
    assign rx_pin[58] = mb1_BA1_IO_046_mb1_BC1_IO_044;

    assign mb1_BA1_IO_047_mb1_BC1_IO_045 = tx_pin[0];
    assign mb1_BA1_IO_048_mb1_BC1_IO_062 = tx_pin[1];
    assign mb1_BA1_IO_049_mb1_BC1_IO_063 = tx_pin[2];
    assign mb1_BA1_IO_050_mb1_BC1_IO_040 = tx_pin[3];
    assign mb1_BA1_IO_051_mb1_BC1_IO_041 = tx_pin[4];
    assign mb1_BA1_IO_052_mb1_BC1_IO_038 = tx_pin[5];
    assign mb1_BA1_IO_053_mb1_BC1_IO_039 = tx_pin[6];
    assign mb1_BA1_IO_054_mb1_BC1_IO_056 = tx_pin[7];
    assign mb1_BA1_IO_055_mb1_BC1_IO_057 = tx_pin[8];
    assign mb1_BA1_IO_056_mb1_BC1_IO_054 = tx_pin[9];
    assign mb1_BA1_IO_057_mb1_BC1_IO_055 = tx_pin[10];
    assign mb1_BA1_IO_058_mb1_BC1_IO_072 = tx_pin[11];
    assign mb1_BA1_IO_059_mb1_BC1_IO_073 = tx_pin[12];
    assign mb1_BA1_IO_060_mb1_BC1_IO_070 = tx_pin[13];
    assign mb1_BA1_IO_061_mb1_BC1_IO_071 = tx_pin[14];
    assign mb1_BA1_IO_062_mb1_BC1_IO_048 = tx_pin[15];
    assign mb1_BA1_IO_063_mb1_BC1_IO_049 = tx_pin[16];
    assign mb1_BA1_IO_064_mb1_BC1_IO_066 = tx_pin[17];
    assign mb1_BA1_IO_065_mb1_BC1_IO_067 = tx_pin[18];
    assign mb1_BA1_IO_066_mb1_BC1_IO_064 = tx_pin[19];
    assign mb1_BA1_IO_067_mb1_BC1_IO_065 = tx_pin[20];
    assign mb1_BA1_IO_068_mb1_BC1_IO_082 = tx_pin[21];
    assign mb1_BA1_IO_069_mb1_BC1_IO_083 = tx_pin[22];
    assign mb1_BA1_IO_070_mb1_BC1_IO_060 = tx_pin[23];
    assign mb1_BA1_IO_071_mb1_BC1_IO_061 = tx_pin[24];
    assign mb1_BA1_IO_072_mb1_BC1_IO_058 = tx_pin[25];
    assign mb1_BA1_IO_073_mb1_BC1_IO_059 = tx_pin[26];
    assign mb1_BA1_IO_074_mb1_BC1_IO_076 = tx_pin[27];
    assign mb1_BA1_IO_075_mb1_BC1_IO_077 = tx_pin[28];
    assign mb1_BA1_IO_076_mb1_BC1_IO_074 = tx_pin[29];
    assign mb1_BA1_IO_077_mb1_BC1_IO_075 = tx_pin[30];
    assign mb1_BA1_IO_078_mb1_BC1_IO_092 = tx_pin[31];
    assign mb1_BA1_IO_079_mb1_BC1_IO_093 = tx_pin[32];
    assign mb1_BA1_IO_080_mb1_BC1_IO_090 = tx_pin[33];
    assign mb1_BA1_IO_081_mb1_BC1_IO_091 = tx_pin[34];
    assign mb1_BA1_IO_082_mb1_BC1_IO_068 = tx_pin[35];
    assign mb1_BA1_IO_083_mb1_BC1_IO_069 = tx_pin[36];
    assign mb1_BA1_IO_084_mb1_BC1_IO_086 = tx_pin[37];
    assign mb1_BA1_IO_085_mb1_BC1_IO_087 = tx_pin[38];
    assign mb1_BA1_IO_086_mb1_BC1_IO_084 = tx_pin[39];
    assign mb1_BA1_IO_087_mb1_BC1_IO_085 = tx_pin[40];
    assign mb1_BA1_IO_088_mb1_BC1_IO_102 = tx_pin[41];
    assign mb1_BA1_IO_089_mb1_BC1_IO_103 = tx_pin[42];
    assign mb1_BA1_IO_090_mb1_BC1_IO_080 = tx_pin[43];
    assign mb1_BA1_IO_091_mb1_BC1_IO_081 = tx_pin[44];
    assign mb1_BA1_IO_092_mb1_BC1_IO_078 = tx_pin[45];
    assign mb1_BA1_IO_093_mb1_BC1_IO_079 = tx_pin[46];
    assign mb1_BA1_IO_094_mb1_BC1_IO_096 = tx_pin[47];
    assign mb1_BA1_IO_095_mb1_BC1_IO_097 = tx_pin[48];
    assign mb1_BA1_IO_096_mb1_BC1_IO_094 = tx_pin[49];
    assign mb1_BA1_IO_097_mb1_BC1_IO_095 = tx_pin[50];
    assign mb1_BA1_IO_098_mb1_BC1_IO_112 = tx_pin[51];
    assign mb1_BA1_IO_099_mb1_BC1_IO_113 = tx_pin[52];
    assign mb1_BA1_IO_100_mb1_BC1_IO_110 = tx_pin[53];
    assign mb1_BA1_IO_101_mb1_BC1_IO_111 = tx_pin[54];
    assign mb1_BA1_IO_102_mb1_BC1_IO_088 = tx_pin[55];
    assign mb1_BA1_IO_103_mb1_BC1_IO_089 = tx_pin[56];
    assign mb1_BA1_IO_104_mb1_BC1_IO_106 = tx_pin[57];
    assign mb1_BA1_IO_105_mb1_BC1_IO_107 = tx_pin[58];

    wire [TX_PINS-1:0] tx2_pin;
    wire [RX_PINS-1:0] rx2_pin;

    /* pins which are connected to motherboard connector BB1 */
    /* and connector BA1 on x-board IC-PDS-CABLE-R1 */
    assign rx2_pin[0] = mb1_BB1_CLKIO_N_0_mb1_BB3_CLKIO_N_7;
    assign rx2_pin[1] = mb1_BB1_CLKIO_N_1_mb1_BB3_CLKIO_N_6;
    assign rx2_pin[2] = mb1_BB1_CLKIO_N_2_mb1_BB3_CLKIO_N_4;
    assign rx2_pin[3] = mb1_BB1_CLKIO_N_3_mb1_BB3_CLKIO_N_3;
    assign rx2_pin[4] = mb1_BB1_CLKIO_N_4_mb1_BB3_CLKIO_N_2;
    assign rx2_pin[5] = mb1_BB1_CLKIO_N_5_mb1_BB3_IO_010;
    assign rx2_pin[6] = mb1_BB1_CLKIO_N_6_mb1_BB3_CLKIO_N_1;
    assign rx2_pin[7] = mb1_BB1_CLKIO_N_7_mb1_BB3_CLKIO_N_0;
    assign rx2_pin[8] = mb1_BB1_CLKIO_P_0_mb1_BB3_CLKIO_P_7;
    assign rx2_pin[9] = mb1_BB1_CLKIO_P_1_mb1_BB3_CLKIO_P_6;
    assign rx2_pin[10] = mb1_BB1_CLKIO_P_2_mb1_BB3_CLKIO_P_4;
    assign rx2_pin[11] = mb1_BB1_CLKIO_P_3_mb1_BB3_CLKIO_P_3;
    assign rx2_pin[12] = mb1_BB1_CLKIO_P_4_mb1_BB3_CLKIO_P_2;
    assign rx2_pin[13] = mb1_BB1_CLKIO_P_5_mb1_BB3_IO_011;
    assign rx2_pin[14] = mb1_BB1_CLKIO_P_6_mb1_BB3_CLKIO_P_1;
    assign rx2_pin[15] = mb1_BB1_CLKIO_P_7_mb1_BB3_CLKIO_P_0;
    assign rx2_pin[16] = mb1_BB1_IO_004_mb1_BB3_IO_006;
    assign rx2_pin[17] = mb1_BB1_IO_005_mb1_BB3_IO_007;
    assign rx2_pin[18] = mb1_BB1_IO_006_mb1_BB3_IO_004;
    assign rx2_pin[19] = mb1_BB1_IO_007_mb1_BB3_IO_005;
    assign rx2_pin[20] = mb1_BB1_IO_008_mb1_BB3_IO_022;
    assign rx2_pin[21] = mb1_BB1_IO_009_mb1_BB3_IO_023;
    assign rx2_pin[22] = mb1_BB1_IO_010_mb1_BB3_CLKIO_N_5;
    assign rx2_pin[23] = mb1_BB1_IO_011_mb1_BB3_CLKIO_P_5;
    assign rx2_pin[24] = mb1_BB1_IO_012_mb1_BB3_IO_012;
    assign rx2_pin[25] = mb1_BB1_IO_013_mb1_BB3_IO_013;
    assign rx2_pin[26] = mb1_BB1_IO_014_mb1_BB3_IO_016;
    assign rx2_pin[27] = mb1_BB1_IO_015_mb1_BB3_IO_017;
    assign rx2_pin[28] = mb1_BB1_IO_016_mb1_BB3_IO_014;
    assign rx2_pin[29] = mb1_BB1_IO_017_mb1_BB3_IO_015;
    assign rx2_pin[30] = mb1_BB1_IO_018_mb1_BB3_IO_032;
    assign rx2_pin[31] = mb1_BB1_IO_019_mb1_BB3_IO_033;
    assign rx2_pin[32] = mb1_BB1_IO_020_mb1_BB3_IO_030;
    assign rx2_pin[33] = mb1_BB1_IO_021_mb1_BB3_IO_031;
    assign rx2_pin[34] = mb1_BB1_IO_022_mb1_BB3_IO_008;
    assign rx2_pin[35] = mb1_BB1_IO_023_mb1_BB3_IO_009;
    assign rx2_pin[36] = mb1_BB1_IO_024_mb1_BB3_IO_026;
    assign rx2_pin[37] = mb1_BB1_IO_025_mb1_BB3_IO_027;
    assign rx2_pin[38] = mb1_BB1_IO_026_mb1_BB3_IO_024;
    assign rx2_pin[39] = mb1_BB1_IO_027_mb1_BB3_IO_025;
    assign rx2_pin[40] = mb1_BB1_IO_028_mb1_BB3_IO_042;
    assign rx2_pin[41] = mb1_BB1_IO_029_mb1_BB3_IO_043;
    assign rx2_pin[42] = mb1_BB1_IO_030_mb1_BB3_IO_020;
    assign rx2_pin[43] = mb1_BB1_IO_031_mb1_BB3_IO_021;
    assign rx2_pin[44] = mb1_BB1_IO_032_mb1_BB3_IO_018;
    assign rx2_pin[45] = mb1_BB1_IO_033_mb1_BB3_IO_019;
    assign rx2_pin[46] = mb1_BB1_IO_034_mb1_BB3_IO_036;
    assign rx2_pin[47] = mb1_BB1_IO_035_mb1_BB3_IO_037;
    assign rx2_pin[48] = mb1_BB1_IO_036_mb1_BB3_IO_034;
    assign rx2_pin[49] = mb1_BB1_IO_037_mb1_BB3_IO_035;
    assign rx2_pin[50] = mb1_BB1_IO_038_mb1_BB3_IO_052;
    assign rx2_pin[51] = mb1_BB1_IO_039_mb1_BB3_IO_053;
    assign rx2_pin[52] = mb1_BB1_IO_040_mb1_BB3_IO_050;
    assign rx2_pin[53] = mb1_BB1_IO_041_mb1_BB3_IO_051;
    assign rx2_pin[54] = mb1_BB1_IO_042_mb1_BB3_IO_028;
    assign rx2_pin[55] = mb1_BB1_IO_043_mb1_BB3_IO_029;
    assign rx2_pin[56] = mb1_BB1_IO_044_mb1_BB3_IO_046;
    assign rx2_pin[57] = mb1_BB1_IO_045_mb1_BB3_IO_047;
    assign rx2_pin[58] = mb1_BB1_IO_046_mb1_BB3_IO_044;

    assign mb1_BB1_IO_047_mb1_BB3_IO_045 = tx2_pin[0];
    assign mb1_BB1_IO_048_mb1_BB3_IO_062 = tx2_pin[1];
    assign mb1_BB1_IO_049_mb1_BB3_IO_063 = tx2_pin[2];
    assign mb1_BB1_IO_050_mb1_BB3_IO_040 = tx2_pin[3];
    assign mb1_BB1_IO_051_mb1_BB3_IO_041 = tx2_pin[4];
    assign mb1_BB1_IO_052_mb1_BB3_IO_038 = tx2_pin[5];
    assign mb1_BB1_IO_053_mb1_BB3_IO_039 = tx2_pin[6];
    assign mb1_BB1_IO_054_mb1_BB3_IO_056 = tx2_pin[7];
    assign mb1_BB1_IO_055_mb1_BB3_IO_057 = tx2_pin[8];
    assign mb1_BB1_IO_056_mb1_BB3_IO_054 = tx2_pin[9];
    assign mb1_BB1_IO_057_mb1_BB3_IO_055 = tx2_pin[10];
    assign mb1_BB1_IO_058_mb1_BB3_IO_072 = tx2_pin[11];
    assign mb1_BB1_IO_059_mb1_BB3_IO_073 = tx2_pin[12];
    assign mb1_BB1_IO_060_mb1_BB3_IO_070 = tx2_pin[13];
    assign mb1_BB1_IO_061_mb1_BB3_IO_071 = tx2_pin[14];
    assign mb1_BB1_IO_062_mb1_BB3_IO_048 = tx2_pin[15];
    assign mb1_BB1_IO_063_mb1_BB3_IO_049 = tx2_pin[16];
    assign mb1_BB1_IO_064_mb1_BB3_IO_066 = tx2_pin[17];
    assign mb1_BB1_IO_065_mb1_BB3_IO_067 = tx2_pin[18];
    assign mb1_BB1_IO_066_mb1_BB3_IO_064 = tx2_pin[19];
    assign mb1_BB1_IO_067_mb1_BB3_IO_065 = tx2_pin[20];
    assign mb1_BB1_IO_068_mb1_BB3_IO_082 = tx2_pin[21];
    assign mb1_BB1_IO_069_mb1_BB3_IO_083 = tx2_pin[22];
    assign mb1_BB1_IO_070_mb1_BB3_IO_060 = tx2_pin[23];
    assign mb1_BB1_IO_071_mb1_BB3_IO_061 = tx2_pin[24];
    assign mb1_BB1_IO_072_mb1_BB3_IO_058 = tx2_pin[25];
    assign mb1_BB1_IO_073_mb1_BB3_IO_059 = tx2_pin[26];
    assign mb1_BB1_IO_074_mb1_BB3_IO_076 = tx2_pin[27];
    assign mb1_BB1_IO_075_mb1_BB3_IO_077 = tx2_pin[28];
    assign mb1_BB1_IO_076_mb1_BB3_IO_074 = tx2_pin[29];
    assign mb1_BB1_IO_077_mb1_BB3_IO_075 = tx2_pin[30];
    assign mb1_BB1_IO_078_mb1_BB3_IO_092 = tx2_pin[31];
    assign mb1_BB1_IO_079_mb1_BB3_IO_093 = tx2_pin[32];
    assign mb1_BB1_IO_080_mb1_BB3_IO_090 = tx2_pin[33];
    assign mb1_BB1_IO_081_mb1_BB3_IO_091 = tx2_pin[34];
    assign mb1_BB1_IO_082_mb1_BB3_IO_068 = tx2_pin[35];
    assign mb1_BB1_IO_083_mb1_BB3_IO_069 = tx2_pin[36];
    assign mb1_BB1_IO_084_mb1_BB3_IO_086 = tx2_pin[37];
    assign mb1_BB1_IO_085_mb1_BB3_IO_087 = tx2_pin[38];
    assign mb1_BB1_IO_086_mb1_BB3_IO_084 = tx2_pin[39];
    assign mb1_BB1_IO_087_mb1_BB3_IO_085 = tx2_pin[40];
    assign mb1_BB1_IO_088_mb1_BB3_IO_102 = tx2_pin[41];
    assign mb1_BB1_IO_089_mb1_BB3_IO_103 = tx2_pin[42];
    assign mb1_BB1_IO_090_mb1_BB3_IO_080 = tx2_pin[43];
    assign mb1_BB1_IO_091_mb1_BB3_IO_081 = tx2_pin[44];
    assign mb1_BB1_IO_092_mb1_BB3_IO_078 = tx2_pin[45];
    assign mb1_BB1_IO_093_mb1_BB3_IO_079 = tx2_pin[46];
    assign mb1_BB1_IO_094_mb1_BB3_IO_096 = tx2_pin[47];
    assign mb1_BB1_IO_095_mb1_BB3_IO_097 = tx2_pin[48];
    assign mb1_BB1_IO_096_mb1_BB3_IO_094 = tx2_pin[49];
    assign mb1_BB1_IO_097_mb1_BB3_IO_095 = tx2_pin[50];
    assign mb1_BB1_IO_098_mb1_BB3_IO_112 = tx2_pin[51];
    assign mb1_BB1_IO_099_mb1_BB3_IO_113 = tx2_pin[52];
    assign mb1_BB1_IO_100_mb1_BB3_IO_110 = tx2_pin[53];
    assign mb1_BB1_IO_101_mb1_BB3_IO_111 = tx2_pin[54];
    assign mb1_BB1_IO_102_mb1_BB3_IO_088 = tx2_pin[55];
    assign mb1_BB1_IO_103_mb1_BB3_IO_089 = tx2_pin[56];
    assign mb1_BB1_IO_104_mb1_BB3_IO_106 = tx2_pin[57];
    assign mb1_BB1_IO_105_mb1_BB3_IO_107 = tx2_pin[58];

    top #(
        .FPGA(TA1),
        .fpga_x(1),
        .fpga_y(0))
    top_inst (
        .clk0_p(clk0_p),
        .clk0_n(clk0_n),

        .sync0_p(sync0_p),
        .sync0_n(sync0_n),

        .dmbi_h2f(dmbi_h2f),
        .dmbi_f2h(dmbi_f2h),

        .tx_pin(tx_pin),
        .rx_pin(rx_pin),

        .tx2_pin(tx2_pin),
        .rx2_pin(rx2_pin),

        .clk1_p(clk1_p),
        .clk1_n(clk1_n),

        .sync1_p(sync1_p),
        .sync1_n(sync1_n),

        .led_red(led_red),
        .led_green(led_green),
        .led_blue(led_blue),
        .led_yellow(led_yellow),

        `ifdef EN_DDR
            .clk2_p(clk2_p),
            .clk2_n(clk2_n),
        `endif

        // SSRAM interface
        .sram0_k_p(sram0_k_p),
        .sram0_k_n(sram0_k_n),
        .sram0_a(sram0_a),
        .sram0_dq(sram0_dq),
        .sram0_bws_n(sram0_bws_n),
        .sram0_rnw(sram0_rnw),
        .sram0_ld_n(sram0_ld_n),
        .sram0_doff_n(sram0_doff_n),

        .sram1_k_p(sram1_k_p),
        .sram1_k_n(sram1_k_n),
        .sram1_a(sram1_a),
        .sram1_dq(sram1_dq),
        .sram1_bws_n(sram1_bws_n),
        .sram1_rnw(sram1_rnw),
        .sram1_ld_n(sram1_ld_n),
        .sram1_doff_n(sram1_doff_n),

        .sram2_k_p(sram2_k_p),
        .sram2_k_n(sram2_k_n),
        .sram2_a(sram2_a),
        .sram2_dq(sram2_dq),
        .sram2_bws_n(sram2_bws_n),
        .sram2_rnw(sram2_rnw),
        .sram2_ld_n(sram2_ld_n),
        .sram2_doff_n(sram2_doff_n),

        .sram3_k_p(sram3_k_p),
        .sram3_k_n(sram3_k_n),
        .sram3_a(sram3_a),
        .sram3_dq(sram3_dq),
        .sram3_bws_n(sram3_bws_n),
        .sram3_rnw(sram3_rnw),
        .sram3_ld_n(sram3_ld_n),
        .sram3_doff_n(sram3_doff_n)

        `ifdef EN_DDR
            ,
            .ddr3_dq(ddr3_dq),
            .ddr3_dqs_p(ddr3_dqs_p),
            .ddr3_dqs_n(ddr3_dqs_n),
            .ddr3_addr(ddr3_addr),
            .ddr3_ba(ddr3_ba),
            .ddr3_ras_n(ddr3_ras_n),
            .ddr3_cas_n(ddr3_cas_n),
            .ddr3_we_n(ddr3_we_n),
            .ddr3_reset_n(ddr3_reset_n),
            .ddr3_ck_p(ddr3_ck_p),
            .ddr3_ck_n(ddr3_ck_n),
            .ddr3_cke(ddr3_cke),
            .ddr3_cs_n(ddr3_cs_n),
            .ddr3_dm(ddr3_dm),
            .ddr3_odt(ddr3_odt)
        `endif

        `ifdef EN_ETH
            ,
            .eth_clk_to_mac(eth_clk_to_mac),
            .eth_col_clk_mac_freq(eth_col_clk_mac_freq),
            .eth_crs_rgmii_sel0(eth_crs_rgmii_sel0),
            .eth_gtx_clk_tck(eth_gtx_clk_tck),
            .eth_mdc(eth_mdc),
            .eth_mdio(eth_mdio),
            .eth_ninterrupt(eth_ninterrupt),
            .eth_nreset(eth_nreset),
            .eth_rx_clk(eth_rx_clk),
            .eth_rx_dv_rck(eth_rx_dv_rck),
            .eth_rx_er_rxdv_er(eth_rx_er_rxdv_er),
            .eth_rxd(eth_rxd),
            .eth_tx_clk_rgmii_sel1(eth_tx_clk_rgmii_sel1),
            .eth_tx_en_txen_er(eth_tx_en_txen_er),
            .eth_tx_er(eth_tx_er),
            .eth_txd(eth_txd)
        `endif
    );
endmodule
